compare_12_inst : compare_12 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AgB	 => AgB_sig
	);
