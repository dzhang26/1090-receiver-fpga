shift_reg_112_1_inst : shift_reg_112_1 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		enable	 => enable_sig,
		sclr	 => sclr_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
