-------------------------------------------------------------------
-- This file is designed for the firmware part of 1.09GHz receiver.
-- Design and implement by Dabin Zhang, all rights reserved.
-------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;  -- DO NOT use "std_logic_signed"

-- 12-bit 400-word shift register
entity shift_reg_400_14 is port
(
	clk,reset: in std_logic;
	data_in: in std_logic_vector(13 downto 0);
	-- ,data_376,data_374  -- removed @ 201307272122
	data_399,data_391,data_383,data_375,data_367,data_359: out std_logic_vector(13 downto 0)
);
end shift_reg_400_14;

architecture behavioral of shift_reg_400_14 is

signal reg_399_signal,reg_398_signal,reg_397_signal,reg_396_signal,reg_395_signal,reg_394_signal,reg_393_signal,reg_392_signal,reg_391_signal,reg_390_signal,reg_389_signal,reg_388_signal,reg_387_signal,reg_386_signal,reg_385_signal,reg_384_signal,reg_383_signal,reg_382_signal,reg_381_signal,reg_380_signal,reg_379_signal,reg_378_signal,reg_377_signal,reg_376_signal,reg_375_signal,reg_374_signal,reg_373_signal,reg_372_signal,reg_371_signal,reg_370_signal,reg_369_signal,reg_368_signal,reg_367_signal,reg_366_signal,reg_365_signal,reg_364_signal,reg_363_signal,reg_362_signal,reg_361_signal,reg_360_signal,reg_359_signal,reg_358_signal,reg_357_signal,reg_356_signal,reg_355_signal,reg_354_signal,reg_353_signal,reg_352_signal,reg_351_signal,reg_350_signal,reg_349_signal,reg_348_signal,reg_347_signal,reg_346_signal,reg_345_signal,reg_344_signal,reg_343_signal,reg_342_signal,reg_341_signal,reg_340_signal,reg_339_signal,reg_338_signal,reg_337_signal,reg_336_signal,reg_335_signal,reg_334_signal,reg_333_signal,reg_332_signal,reg_331_signal,reg_330_signal,reg_329_signal,reg_328_signal,reg_327_signal,reg_326_signal,reg_325_signal,reg_324_signal,reg_323_signal,reg_322_signal,reg_321_signal,reg_320_signal,reg_319_signal,reg_318_signal,reg_317_signal,reg_316_signal,reg_315_signal,reg_314_signal,reg_313_signal,reg_312_signal,reg_311_signal,reg_310_signal,reg_309_signal,reg_308_signal,reg_307_signal,reg_306_signal,reg_305_signal,reg_304_signal,reg_303_signal,reg_302_signal,reg_301_signal,reg_300_signal,
reg_299_signal,reg_298_signal,reg_297_signal,reg_296_signal,reg_295_signal,reg_294_signal,reg_293_signal,reg_292_signal,reg_291_signal,reg_290_signal,reg_289_signal,reg_288_signal,reg_287_signal,reg_286_signal,reg_285_signal,reg_284_signal,reg_283_signal,reg_282_signal,reg_281_signal,reg_280_signal,reg_279_signal,reg_278_signal,reg_277_signal,reg_276_signal,reg_275_signal,reg_274_signal,reg_273_signal,reg_272_signal,reg_271_signal,reg_270_signal,reg_269_signal,reg_268_signal,reg_267_signal,reg_266_signal,reg_265_signal,reg_264_signal,reg_263_signal,reg_262_signal,reg_261_signal,reg_260_signal,reg_259_signal,reg_258_signal,reg_257_signal,reg_256_signal,reg_255_signal,reg_254_signal,reg_253_signal,reg_252_signal,reg_251_signal,reg_250_signal,reg_249_signal,reg_248_signal,reg_247_signal,reg_246_signal,reg_245_signal,reg_244_signal,reg_243_signal,reg_242_signal,reg_241_signal,reg_240_signal,reg_239_signal,reg_238_signal,reg_237_signal,reg_236_signal,reg_235_signal,reg_234_signal,reg_233_signal,reg_232_signal,reg_231_signal,reg_230_signal,reg_229_signal,reg_228_signal,reg_227_signal,reg_226_signal,reg_225_signal,reg_224_signal,reg_223_signal,reg_222_signal,reg_221_signal,reg_220_signal,reg_219_signal,reg_218_signal,reg_217_signal,reg_216_signal,reg_215_signal,reg_214_signal,reg_213_signal,reg_212_signal,reg_211_signal,reg_210_signal,reg_209_signal,reg_208_signal,reg_207_signal,reg_206_signal,reg_205_signal,reg_204_signal,reg_203_signal,reg_202_signal,reg_201_signal,reg_200_signal,
reg_199_signal,reg_198_signal,reg_197_signal,reg_196_signal,reg_195_signal,reg_194_signal,reg_193_signal,reg_192_signal,reg_191_signal,reg_190_signal,reg_189_signal,reg_188_signal,reg_187_signal,reg_186_signal,reg_185_signal,reg_184_signal,reg_183_signal,reg_182_signal,reg_181_signal,reg_180_signal,reg_179_signal,reg_178_signal,reg_177_signal,reg_176_signal,reg_175_signal,reg_174_signal,reg_173_signal,reg_172_signal,reg_171_signal,reg_170_signal,reg_169_signal,reg_168_signal,reg_167_signal,reg_166_signal,reg_165_signal,reg_164_signal,reg_163_signal,reg_162_signal,reg_161_signal,reg_160_signal,reg_159_signal,reg_158_signal,reg_157_signal,reg_156_signal,reg_155_signal,reg_154_signal,reg_153_signal,reg_152_signal,reg_151_signal,reg_150_signal,reg_149_signal,reg_148_signal,reg_147_signal,reg_146_signal,reg_145_signal,reg_144_signal,reg_143_signal,reg_142_signal,reg_141_signal,reg_140_signal,reg_139_signal,reg_138_signal,reg_137_signal,reg_136_signal,reg_135_signal,reg_134_signal,reg_133_signal,reg_132_signal,reg_131_signal,reg_130_signal,reg_129_signal,reg_128_signal,reg_127_signal,reg_126_signal,reg_125_signal,reg_124_signal,reg_123_signal,reg_122_signal,reg_121_signal,reg_120_signal,reg_119_signal,reg_118_signal,reg_117_signal,reg_116_signal,reg_115_signal,reg_114_signal,reg_113_signal,reg_112_signal,reg_111_signal,reg_110_signal,reg_109_signal,reg_108_signal,reg_107_signal,reg_106_signal,reg_105_signal,reg_104_signal,reg_103_signal,reg_102_signal,reg_101_signal,reg_100_signal,
reg_99_signal,reg_98_signal,reg_97_signal,reg_96_signal,reg_95_signal,reg_94_signal,reg_93_signal,reg_92_signal,reg_91_signal,reg_90_signal,reg_89_signal,reg_88_signal,reg_87_signal,reg_86_signal,reg_85_signal,reg_84_signal,reg_83_signal,reg_82_signal,reg_81_signal,reg_80_signal,reg_79_signal,reg_78_signal,reg_77_signal,reg_76_signal,reg_75_signal,reg_74_signal,reg_73_signal,reg_72_signal,reg_71_signal,reg_70_signal,reg_69_signal,reg_68_signal,reg_67_signal,reg_66_signal,reg_65_signal,reg_64_signal,reg_63_signal,reg_62_signal,reg_61_signal,reg_60_signal,reg_59_signal,reg_58_signal,reg_57_signal,reg_56_signal,reg_55_signal,reg_54_signal,reg_53_signal,reg_52_signal,reg_51_signal,reg_50_signal,reg_49_signal,reg_48_signal,reg_47_signal,reg_46_signal,reg_45_signal,reg_44_signal,reg_43_signal,reg_42_signal,reg_41_signal,reg_40_signal,reg_39_signal,reg_38_signal,reg_37_signal,reg_36_signal,reg_35_signal,reg_34_signal,reg_33_signal,reg_32_signal,reg_31_signal,reg_30_signal,reg_29_signal,reg_28_signal,reg_27_signal,reg_26_signal,reg_25_signal,reg_24_signal,reg_23_signal,reg_22_signal,reg_21_signal,reg_20_signal,reg_19_signal,reg_18_signal,reg_17_signal,reg_16_signal,reg_15_signal,reg_14_signal,reg_13_signal,reg_12_signal,reg_11_signal,reg_10_signal,reg_9_signal,reg_8_signal,reg_7_signal,reg_6_signal,reg_5_signal,reg_4_signal,reg_3_signal,reg_2_signal,reg_1_signal,reg_0_signal: std_logic_vector(13 downto 0);

component dff_14 is port
(
	aclr: in std_logic;
	clock: in std_logic;
	data: in std_logic_vector(13 downto 0);
	q: out std_logic_vector(13 downto 0)
);
end component;

begin

reg_399: dff_14 port map(aclr=>reset,clock=>clk,data=>data_in,q=>reg_399_signal);
reg_398: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_399_signal,q=>reg_398_signal);
reg_397: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_398_signal,q=>reg_397_signal);
reg_396: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_397_signal,q=>reg_396_signal);
reg_395: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_396_signal,q=>reg_395_signal);
reg_394: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_395_signal,q=>reg_394_signal);
reg_393: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_394_signal,q=>reg_393_signal);
reg_392: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_393_signal,q=>reg_392_signal);
reg_391: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_392_signal,q=>reg_391_signal);
reg_390: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_391_signal,q=>reg_390_signal);
reg_389: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_390_signal,q=>reg_389_signal);
reg_388: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_389_signal,q=>reg_388_signal);
reg_387: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_388_signal,q=>reg_387_signal);
reg_386: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_387_signal,q=>reg_386_signal);
reg_385: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_386_signal,q=>reg_385_signal);
reg_384: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_385_signal,q=>reg_384_signal);
reg_383: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_384_signal,q=>reg_383_signal);
reg_382: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_383_signal,q=>reg_382_signal);
reg_381: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_382_signal,q=>reg_381_signal);
reg_380: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_381_signal,q=>reg_380_signal);
reg_379: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_380_signal,q=>reg_379_signal);
reg_378: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_379_signal,q=>reg_378_signal);
reg_377: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_378_signal,q=>reg_377_signal);
reg_376: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_377_signal,q=>reg_376_signal);
reg_375: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_376_signal,q=>reg_375_signal);
reg_374: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_375_signal,q=>reg_374_signal);
reg_373: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_374_signal,q=>reg_373_signal);
reg_372: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_373_signal,q=>reg_372_signal);
reg_371: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_372_signal,q=>reg_371_signal);
reg_370: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_371_signal,q=>reg_370_signal);
reg_369: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_370_signal,q=>reg_369_signal);
reg_368: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_369_signal,q=>reg_368_signal);
reg_367: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_368_signal,q=>reg_367_signal);
reg_366: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_367_signal,q=>reg_366_signal);
reg_365: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_366_signal,q=>reg_365_signal);
reg_364: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_365_signal,q=>reg_364_signal);
reg_363: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_364_signal,q=>reg_363_signal);
reg_362: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_363_signal,q=>reg_362_signal);
reg_361: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_362_signal,q=>reg_361_signal);
reg_360: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_361_signal,q=>reg_360_signal);
reg_359: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_360_signal,q=>reg_359_signal);
reg_358: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_359_signal,q=>reg_358_signal);
reg_357: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_358_signal,q=>reg_357_signal);
reg_356: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_357_signal,q=>reg_356_signal);
reg_355: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_356_signal,q=>reg_355_signal);
reg_354: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_355_signal,q=>reg_354_signal);
reg_353: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_354_signal,q=>reg_353_signal);
reg_352: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_353_signal,q=>reg_352_signal);
reg_351: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_352_signal,q=>reg_351_signal);
reg_350: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_351_signal,q=>reg_350_signal);
reg_349: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_350_signal,q=>reg_349_signal);
reg_348: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_349_signal,q=>reg_348_signal);
reg_347: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_348_signal,q=>reg_347_signal);
reg_346: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_347_signal,q=>reg_346_signal);
reg_345: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_346_signal,q=>reg_345_signal);
reg_344: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_345_signal,q=>reg_344_signal);
reg_343: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_344_signal,q=>reg_343_signal);
reg_342: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_343_signal,q=>reg_342_signal);
reg_341: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_342_signal,q=>reg_341_signal);
reg_340: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_341_signal,q=>reg_340_signal);
reg_339: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_340_signal,q=>reg_339_signal);
reg_338: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_339_signal,q=>reg_338_signal);
reg_337: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_338_signal,q=>reg_337_signal);
reg_336: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_337_signal,q=>reg_336_signal);
reg_335: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_336_signal,q=>reg_335_signal);
reg_334: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_335_signal,q=>reg_334_signal);
reg_333: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_334_signal,q=>reg_333_signal);
reg_332: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_333_signal,q=>reg_332_signal);
reg_331: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_332_signal,q=>reg_331_signal);
reg_330: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_331_signal,q=>reg_330_signal);
reg_329: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_330_signal,q=>reg_329_signal);
reg_328: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_329_signal,q=>reg_328_signal);
reg_327: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_328_signal,q=>reg_327_signal);
reg_326: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_327_signal,q=>reg_326_signal);
reg_325: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_326_signal,q=>reg_325_signal);
reg_324: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_325_signal,q=>reg_324_signal);
reg_323: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_324_signal,q=>reg_323_signal);
reg_322: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_323_signal,q=>reg_322_signal);
reg_321: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_322_signal,q=>reg_321_signal);
reg_320: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_321_signal,q=>reg_320_signal);
reg_319: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_320_signal,q=>reg_319_signal);
reg_318: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_319_signal,q=>reg_318_signal);
reg_317: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_318_signal,q=>reg_317_signal);
reg_316: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_317_signal,q=>reg_316_signal);
reg_315: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_316_signal,q=>reg_315_signal);
reg_314: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_315_signal,q=>reg_314_signal);
reg_313: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_314_signal,q=>reg_313_signal);
reg_312: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_313_signal,q=>reg_312_signal);
reg_311: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_312_signal,q=>reg_311_signal);
reg_310: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_311_signal,q=>reg_310_signal);
reg_309: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_310_signal,q=>reg_309_signal);
reg_308: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_309_signal,q=>reg_308_signal);
reg_307: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_308_signal,q=>reg_307_signal);
reg_306: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_307_signal,q=>reg_306_signal);
reg_305: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_306_signal,q=>reg_305_signal);
reg_304: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_305_signal,q=>reg_304_signal);
reg_303: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_304_signal,q=>reg_303_signal);
reg_302: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_303_signal,q=>reg_302_signal);
reg_301: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_302_signal,q=>reg_301_signal);
reg_300: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_301_signal,q=>reg_300_signal);
reg_299: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_300_signal,q=>reg_299_signal);
reg_298: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_299_signal,q=>reg_298_signal);
reg_297: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_298_signal,q=>reg_297_signal);
reg_296: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_297_signal,q=>reg_296_signal);
reg_295: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_296_signal,q=>reg_295_signal);
reg_294: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_295_signal,q=>reg_294_signal);
reg_293: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_294_signal,q=>reg_293_signal);
reg_292: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_293_signal,q=>reg_292_signal);
reg_291: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_292_signal,q=>reg_291_signal);
reg_290: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_291_signal,q=>reg_290_signal);
reg_289: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_290_signal,q=>reg_289_signal);
reg_288: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_289_signal,q=>reg_288_signal);
reg_287: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_288_signal,q=>reg_287_signal);
reg_286: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_287_signal,q=>reg_286_signal);
reg_285: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_286_signal,q=>reg_285_signal);
reg_284: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_285_signal,q=>reg_284_signal);
reg_283: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_284_signal,q=>reg_283_signal);
reg_282: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_283_signal,q=>reg_282_signal);
reg_281: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_282_signal,q=>reg_281_signal);
reg_280: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_281_signal,q=>reg_280_signal);
reg_279: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_280_signal,q=>reg_279_signal);
reg_278: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_279_signal,q=>reg_278_signal);
reg_277: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_278_signal,q=>reg_277_signal);
reg_276: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_277_signal,q=>reg_276_signal);
reg_275: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_276_signal,q=>reg_275_signal);
reg_274: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_275_signal,q=>reg_274_signal);
reg_273: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_274_signal,q=>reg_273_signal);
reg_272: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_273_signal,q=>reg_272_signal);
reg_271: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_272_signal,q=>reg_271_signal);
reg_270: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_271_signal,q=>reg_270_signal);
reg_269: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_270_signal,q=>reg_269_signal);
reg_268: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_269_signal,q=>reg_268_signal);
reg_267: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_268_signal,q=>reg_267_signal);
reg_266: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_267_signal,q=>reg_266_signal);
reg_265: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_266_signal,q=>reg_265_signal);
reg_264: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_265_signal,q=>reg_264_signal);
reg_263: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_264_signal,q=>reg_263_signal);
reg_262: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_263_signal,q=>reg_262_signal);
reg_261: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_262_signal,q=>reg_261_signal);
reg_260: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_261_signal,q=>reg_260_signal);
reg_259: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_260_signal,q=>reg_259_signal);
reg_258: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_259_signal,q=>reg_258_signal);
reg_257: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_258_signal,q=>reg_257_signal);
reg_256: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_257_signal,q=>reg_256_signal);
reg_255: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_256_signal,q=>reg_255_signal);
reg_254: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_255_signal,q=>reg_254_signal);
reg_253: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_254_signal,q=>reg_253_signal);
reg_252: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_253_signal,q=>reg_252_signal);
reg_251: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_252_signal,q=>reg_251_signal);
reg_250: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_251_signal,q=>reg_250_signal);
reg_249: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_250_signal,q=>reg_249_signal);
reg_248: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_249_signal,q=>reg_248_signal);
reg_247: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_248_signal,q=>reg_247_signal);
reg_246: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_247_signal,q=>reg_246_signal);
reg_245: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_246_signal,q=>reg_245_signal);
reg_244: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_245_signal,q=>reg_244_signal);
reg_243: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_244_signal,q=>reg_243_signal);
reg_242: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_243_signal,q=>reg_242_signal);
reg_241: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_242_signal,q=>reg_241_signal);
reg_240: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_241_signal,q=>reg_240_signal);
reg_239: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_240_signal,q=>reg_239_signal);
reg_238: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_239_signal,q=>reg_238_signal);
reg_237: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_238_signal,q=>reg_237_signal);
reg_236: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_237_signal,q=>reg_236_signal);
reg_235: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_236_signal,q=>reg_235_signal);
reg_234: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_235_signal,q=>reg_234_signal);
reg_233: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_234_signal,q=>reg_233_signal);
reg_232: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_233_signal,q=>reg_232_signal);
reg_231: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_232_signal,q=>reg_231_signal);
reg_230: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_231_signal,q=>reg_230_signal);
reg_229: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_230_signal,q=>reg_229_signal);
reg_228: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_229_signal,q=>reg_228_signal);
reg_227: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_228_signal,q=>reg_227_signal);
reg_226: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_227_signal,q=>reg_226_signal);
reg_225: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_226_signal,q=>reg_225_signal);
reg_224: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_225_signal,q=>reg_224_signal);
reg_223: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_224_signal,q=>reg_223_signal);
reg_222: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_223_signal,q=>reg_222_signal);
reg_221: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_222_signal,q=>reg_221_signal);
reg_220: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_221_signal,q=>reg_220_signal);
reg_219: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_220_signal,q=>reg_219_signal);
reg_218: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_219_signal,q=>reg_218_signal);
reg_217: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_218_signal,q=>reg_217_signal);
reg_216: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_217_signal,q=>reg_216_signal);
reg_215: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_216_signal,q=>reg_215_signal);
reg_214: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_215_signal,q=>reg_214_signal);
reg_213: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_214_signal,q=>reg_213_signal);
reg_212: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_213_signal,q=>reg_212_signal);
reg_211: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_212_signal,q=>reg_211_signal);
reg_210: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_211_signal,q=>reg_210_signal);
reg_209: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_210_signal,q=>reg_209_signal);
reg_208: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_209_signal,q=>reg_208_signal);
reg_207: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_208_signal,q=>reg_207_signal);
reg_206: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_207_signal,q=>reg_206_signal);
reg_205: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_206_signal,q=>reg_205_signal);
reg_204: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_205_signal,q=>reg_204_signal);
reg_203: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_204_signal,q=>reg_203_signal);
reg_202: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_203_signal,q=>reg_202_signal);
reg_201: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_202_signal,q=>reg_201_signal);
reg_200: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_201_signal,q=>reg_200_signal);
reg_199: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_200_signal,q=>reg_199_signal);
reg_198: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_199_signal,q=>reg_198_signal);
reg_197: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_198_signal,q=>reg_197_signal);
reg_196: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_197_signal,q=>reg_196_signal);
reg_195: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_196_signal,q=>reg_195_signal);
reg_194: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_195_signal,q=>reg_194_signal);
reg_193: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_194_signal,q=>reg_193_signal);
reg_192: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_193_signal,q=>reg_192_signal);
reg_191: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_192_signal,q=>reg_191_signal);
reg_190: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_191_signal,q=>reg_190_signal);
reg_189: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_190_signal,q=>reg_189_signal);
reg_188: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_189_signal,q=>reg_188_signal);
reg_187: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_188_signal,q=>reg_187_signal);
reg_186: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_187_signal,q=>reg_186_signal);
reg_185: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_186_signal,q=>reg_185_signal);
reg_184: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_185_signal,q=>reg_184_signal);
reg_183: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_184_signal,q=>reg_183_signal);
reg_182: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_183_signal,q=>reg_182_signal);
reg_181: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_182_signal,q=>reg_181_signal);
reg_180: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_181_signal,q=>reg_180_signal);
reg_179: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_180_signal,q=>reg_179_signal);
reg_178: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_179_signal,q=>reg_178_signal);
reg_177: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_178_signal,q=>reg_177_signal);
reg_176: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_177_signal,q=>reg_176_signal);
reg_175: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_176_signal,q=>reg_175_signal);
reg_174: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_175_signal,q=>reg_174_signal);
reg_173: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_174_signal,q=>reg_173_signal);
reg_172: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_173_signal,q=>reg_172_signal);
reg_171: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_172_signal,q=>reg_171_signal);
reg_170: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_171_signal,q=>reg_170_signal);
reg_169: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_170_signal,q=>reg_169_signal);
reg_168: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_169_signal,q=>reg_168_signal);
reg_167: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_168_signal,q=>reg_167_signal);
reg_166: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_167_signal,q=>reg_166_signal);
reg_165: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_166_signal,q=>reg_165_signal);
reg_164: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_165_signal,q=>reg_164_signal);
reg_163: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_164_signal,q=>reg_163_signal);
reg_162: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_163_signal,q=>reg_162_signal);
reg_161: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_162_signal,q=>reg_161_signal);
reg_160: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_161_signal,q=>reg_160_signal);
reg_159: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_160_signal,q=>reg_159_signal);
reg_158: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_159_signal,q=>reg_158_signal);
reg_157: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_158_signal,q=>reg_157_signal);
reg_156: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_157_signal,q=>reg_156_signal);
reg_155: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_156_signal,q=>reg_155_signal);
reg_154: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_155_signal,q=>reg_154_signal);
reg_153: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_154_signal,q=>reg_153_signal);
reg_152: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_153_signal,q=>reg_152_signal);
reg_151: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_152_signal,q=>reg_151_signal);
reg_150: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_151_signal,q=>reg_150_signal);
reg_149: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_150_signal,q=>reg_149_signal);
reg_148: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_149_signal,q=>reg_148_signal);
reg_147: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_148_signal,q=>reg_147_signal);
reg_146: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_147_signal,q=>reg_146_signal);
reg_145: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_146_signal,q=>reg_145_signal);
reg_144: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_145_signal,q=>reg_144_signal);
reg_143: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_144_signal,q=>reg_143_signal);
reg_142: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_143_signal,q=>reg_142_signal);
reg_141: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_142_signal,q=>reg_141_signal);
reg_140: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_141_signal,q=>reg_140_signal);
reg_139: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_140_signal,q=>reg_139_signal);
reg_138: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_139_signal,q=>reg_138_signal);
reg_137: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_138_signal,q=>reg_137_signal);
reg_136: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_137_signal,q=>reg_136_signal);
reg_135: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_136_signal,q=>reg_135_signal);
reg_134: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_135_signal,q=>reg_134_signal);
reg_133: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_134_signal,q=>reg_133_signal);
reg_132: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_133_signal,q=>reg_132_signal);
reg_131: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_132_signal,q=>reg_131_signal);
reg_130: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_131_signal,q=>reg_130_signal);
reg_129: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_130_signal,q=>reg_129_signal);
reg_128: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_129_signal,q=>reg_128_signal);
reg_127: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_128_signal,q=>reg_127_signal);
reg_126: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_127_signal,q=>reg_126_signal);
reg_125: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_126_signal,q=>reg_125_signal);
reg_124: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_125_signal,q=>reg_124_signal);
reg_123: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_124_signal,q=>reg_123_signal);
reg_122: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_123_signal,q=>reg_122_signal);
reg_121: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_122_signal,q=>reg_121_signal);
reg_120: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_121_signal,q=>reg_120_signal);
reg_119: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_120_signal,q=>reg_119_signal);
reg_118: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_119_signal,q=>reg_118_signal);
reg_117: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_118_signal,q=>reg_117_signal);
reg_116: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_117_signal,q=>reg_116_signal);
reg_115: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_116_signal,q=>reg_115_signal);
reg_114: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_115_signal,q=>reg_114_signal);
reg_113: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_114_signal,q=>reg_113_signal);
reg_112: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_113_signal,q=>reg_112_signal);
reg_111: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_112_signal,q=>reg_111_signal);
reg_110: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_111_signal,q=>reg_110_signal);
reg_109: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_110_signal,q=>reg_109_signal);
reg_108: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_109_signal,q=>reg_108_signal);
reg_107: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_108_signal,q=>reg_107_signal);
reg_106: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_107_signal,q=>reg_106_signal);
reg_105: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_106_signal,q=>reg_105_signal);
reg_104: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_105_signal,q=>reg_104_signal);
reg_103: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_104_signal,q=>reg_103_signal);
reg_102: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_103_signal,q=>reg_102_signal);
reg_101: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_102_signal,q=>reg_101_signal);
reg_100: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_101_signal,q=>reg_100_signal);
reg_99: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_100_signal,q=>reg_99_signal);
reg_98: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_99_signal,q=>reg_98_signal);
reg_97: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_98_signal,q=>reg_97_signal);
reg_96: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_97_signal,q=>reg_96_signal);
reg_95: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_96_signal,q=>reg_95_signal);
reg_94: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_95_signal,q=>reg_94_signal);
reg_93: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_94_signal,q=>reg_93_signal);
reg_92: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_93_signal,q=>reg_92_signal);
reg_91: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_92_signal,q=>reg_91_signal);
reg_90: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_91_signal,q=>reg_90_signal);
reg_89: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_90_signal,q=>reg_89_signal);
reg_88: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_89_signal,q=>reg_88_signal);
reg_87: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_88_signal,q=>reg_87_signal);
reg_86: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_87_signal,q=>reg_86_signal);
reg_85: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_86_signal,q=>reg_85_signal);
reg_84: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_85_signal,q=>reg_84_signal);
reg_83: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_84_signal,q=>reg_83_signal);
reg_82: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_83_signal,q=>reg_82_signal);
reg_81: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_82_signal,q=>reg_81_signal);
reg_80: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_81_signal,q=>reg_80_signal);
reg_79: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_80_signal,q=>reg_79_signal);
reg_78: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_79_signal,q=>reg_78_signal);
reg_77: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_78_signal,q=>reg_77_signal);
reg_76: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_77_signal,q=>reg_76_signal);
reg_75: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_76_signal,q=>reg_75_signal);
reg_74: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_75_signal,q=>reg_74_signal);
reg_73: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_74_signal,q=>reg_73_signal);
reg_72: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_73_signal,q=>reg_72_signal);
reg_71: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_72_signal,q=>reg_71_signal);
reg_70: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_71_signal,q=>reg_70_signal);
reg_69: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_70_signal,q=>reg_69_signal);
reg_68: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_69_signal,q=>reg_68_signal);
reg_67: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_68_signal,q=>reg_67_signal);
reg_66: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_67_signal,q=>reg_66_signal);
reg_65: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_66_signal,q=>reg_65_signal);
reg_64: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_65_signal,q=>reg_64_signal);
reg_63: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_64_signal,q=>reg_63_signal);
reg_62: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_63_signal,q=>reg_62_signal);
reg_61: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_62_signal,q=>reg_61_signal);
reg_60: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_61_signal,q=>reg_60_signal);
reg_59: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_60_signal,q=>reg_59_signal);
reg_58: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_59_signal,q=>reg_58_signal);
reg_57: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_58_signal,q=>reg_57_signal);
reg_56: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_57_signal,q=>reg_56_signal);
reg_55: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_56_signal,q=>reg_55_signal);
reg_54: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_55_signal,q=>reg_54_signal);
reg_53: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_54_signal,q=>reg_53_signal);
reg_52: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_53_signal,q=>reg_52_signal);
reg_51: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_52_signal,q=>reg_51_signal);
reg_50: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_51_signal,q=>reg_50_signal);
reg_49: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_50_signal,q=>reg_49_signal);
reg_48: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_49_signal,q=>reg_48_signal);
reg_47: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_48_signal,q=>reg_47_signal);
reg_46: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_47_signal,q=>reg_46_signal);
reg_45: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_46_signal,q=>reg_45_signal);
reg_44: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_45_signal,q=>reg_44_signal);
reg_43: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_44_signal,q=>reg_43_signal);
reg_42: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_43_signal,q=>reg_42_signal);
reg_41: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_42_signal,q=>reg_41_signal);
reg_40: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_41_signal,q=>reg_40_signal);
reg_39: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_40_signal,q=>reg_39_signal);
reg_38: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_39_signal,q=>reg_38_signal);
reg_37: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_38_signal,q=>reg_37_signal);
reg_36: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_37_signal,q=>reg_36_signal);
reg_35: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_36_signal,q=>reg_35_signal);
reg_34: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_35_signal,q=>reg_34_signal);
reg_33: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_34_signal,q=>reg_33_signal);
reg_32: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_33_signal,q=>reg_32_signal);
reg_31: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_32_signal,q=>reg_31_signal);
reg_30: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_31_signal,q=>reg_30_signal);
reg_29: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_30_signal,q=>reg_29_signal);
reg_28: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_29_signal,q=>reg_28_signal);
reg_27: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_28_signal,q=>reg_27_signal);
reg_26: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_27_signal,q=>reg_26_signal);
reg_25: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_26_signal,q=>reg_25_signal);
reg_24: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_25_signal,q=>reg_24_signal);
reg_23: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_24_signal,q=>reg_23_signal);
reg_22: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_23_signal,q=>reg_22_signal);
reg_21: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_22_signal,q=>reg_21_signal);
reg_20: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_21_signal,q=>reg_20_signal);
reg_19: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_20_signal,q=>reg_19_signal);
reg_18: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_19_signal,q=>reg_18_signal);
reg_17: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_18_signal,q=>reg_17_signal);
reg_16: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_17_signal,q=>reg_16_signal);
reg_15: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_16_signal,q=>reg_15_signal);
reg_14: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_15_signal,q=>reg_14_signal);
reg_13: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_14_signal,q=>reg_13_signal);
reg_12: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_13_signal,q=>reg_12_signal);
reg_11: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_12_signal,q=>reg_11_signal);
reg_10: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_11_signal,q=>reg_10_signal);
reg_9: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_10_signal,q=>reg_9_signal);
reg_8: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_9_signal,q=>reg_8_signal);
reg_7: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_8_signal,q=>reg_7_signal);
reg_6: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_7_signal,q=>reg_6_signal);
reg_5: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_6_signal,q=>reg_5_signal);
reg_4: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_5_signal,q=>reg_4_signal);
reg_3: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_4_signal,q=>reg_3_signal);
reg_2: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_3_signal,q=>reg_2_signal);
reg_1: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_2_signal,q=>reg_1_signal);
reg_0: dff_14 port map(aclr=>reset,clock=>clk,data=>reg_1_signal,q=>reg_0_signal);

data_399<=reg_399_signal;  --399
data_391<=reg_391_signal;  --391
data_383<=reg_383_signal;  --383
--data_376<=reg_376_signal;  --376
data_375<=reg_375_signal;  --375
--data_374<=reg_374_signal;  --374
data_367<=reg_367_signal;
data_359<=reg_359_signal;

end behavioral;