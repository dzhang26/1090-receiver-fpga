clkctrl_50_inst : clkctrl_50 PORT MAP (
		ena	 => ena_sig,
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
