compare_sign_12_inst : compare_sign_12 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		AgB	 => AgB_sig
	);
