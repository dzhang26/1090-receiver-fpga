mux_51_180_p1_inst : mux_51_180_p1 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		data2x	 => data2x_sig,
		data3x	 => data3x_sig,
		data4x	 => data4x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
