adder_12_inst : adder_12 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
