dff_12_inst : dff_12 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
