reg_24_inst : reg_24 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
