-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: mux_51_180_p1.vhd
-- Megafunction Name(s):
-- 			lpm_mux
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux_51_180_p1 IS
	PORT
	(
		aclr		: IN STD_LOGIC  := '0';
		clock		: IN STD_LOGIC ;
		data0x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (179 DOWNTO 0)
	);
END mux_51_180_p1;


ARCHITECTURE SYN OF mux_51_180_p1 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (4 DOWNTO 0, 179 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (179 DOWNTO 0);

BEGIN
	sub_wire6    <= data0x(179 DOWNTO 0);
	sub_wire5    <= data1x(179 DOWNTO 0);
	sub_wire4    <= data2x(179 DOWNTO 0);
	sub_wire3    <= data3x(179 DOWNTO 0);
	result    <= sub_wire0(179 DOWNTO 0);
	sub_wire1    <= data4x(179 DOWNTO 0);
	sub_wire2(4, 0)    <= sub_wire1(0);
	sub_wire2(4, 1)    <= sub_wire1(1);
	sub_wire2(4, 2)    <= sub_wire1(2);
	sub_wire2(4, 3)    <= sub_wire1(3);
	sub_wire2(4, 4)    <= sub_wire1(4);
	sub_wire2(4, 5)    <= sub_wire1(5);
	sub_wire2(4, 6)    <= sub_wire1(6);
	sub_wire2(4, 7)    <= sub_wire1(7);
	sub_wire2(4, 8)    <= sub_wire1(8);
	sub_wire2(4, 9)    <= sub_wire1(9);
	sub_wire2(4, 10)    <= sub_wire1(10);
	sub_wire2(4, 11)    <= sub_wire1(11);
	sub_wire2(4, 12)    <= sub_wire1(12);
	sub_wire2(4, 13)    <= sub_wire1(13);
	sub_wire2(4, 14)    <= sub_wire1(14);
	sub_wire2(4, 15)    <= sub_wire1(15);
	sub_wire2(4, 16)    <= sub_wire1(16);
	sub_wire2(4, 17)    <= sub_wire1(17);
	sub_wire2(4, 18)    <= sub_wire1(18);
	sub_wire2(4, 19)    <= sub_wire1(19);
	sub_wire2(4, 20)    <= sub_wire1(20);
	sub_wire2(4, 21)    <= sub_wire1(21);
	sub_wire2(4, 22)    <= sub_wire1(22);
	sub_wire2(4, 23)    <= sub_wire1(23);
	sub_wire2(4, 24)    <= sub_wire1(24);
	sub_wire2(4, 25)    <= sub_wire1(25);
	sub_wire2(4, 26)    <= sub_wire1(26);
	sub_wire2(4, 27)    <= sub_wire1(27);
	sub_wire2(4, 28)    <= sub_wire1(28);
	sub_wire2(4, 29)    <= sub_wire1(29);
	sub_wire2(4, 30)    <= sub_wire1(30);
	sub_wire2(4, 31)    <= sub_wire1(31);
	sub_wire2(4, 32)    <= sub_wire1(32);
	sub_wire2(4, 33)    <= sub_wire1(33);
	sub_wire2(4, 34)    <= sub_wire1(34);
	sub_wire2(4, 35)    <= sub_wire1(35);
	sub_wire2(4, 36)    <= sub_wire1(36);
	sub_wire2(4, 37)    <= sub_wire1(37);
	sub_wire2(4, 38)    <= sub_wire1(38);
	sub_wire2(4, 39)    <= sub_wire1(39);
	sub_wire2(4, 40)    <= sub_wire1(40);
	sub_wire2(4, 41)    <= sub_wire1(41);
	sub_wire2(4, 42)    <= sub_wire1(42);
	sub_wire2(4, 43)    <= sub_wire1(43);
	sub_wire2(4, 44)    <= sub_wire1(44);
	sub_wire2(4, 45)    <= sub_wire1(45);
	sub_wire2(4, 46)    <= sub_wire1(46);
	sub_wire2(4, 47)    <= sub_wire1(47);
	sub_wire2(4, 48)    <= sub_wire1(48);
	sub_wire2(4, 49)    <= sub_wire1(49);
	sub_wire2(4, 50)    <= sub_wire1(50);
	sub_wire2(4, 51)    <= sub_wire1(51);
	sub_wire2(4, 52)    <= sub_wire1(52);
	sub_wire2(4, 53)    <= sub_wire1(53);
	sub_wire2(4, 54)    <= sub_wire1(54);
	sub_wire2(4, 55)    <= sub_wire1(55);
	sub_wire2(4, 56)    <= sub_wire1(56);
	sub_wire2(4, 57)    <= sub_wire1(57);
	sub_wire2(4, 58)    <= sub_wire1(58);
	sub_wire2(4, 59)    <= sub_wire1(59);
	sub_wire2(4, 60)    <= sub_wire1(60);
	sub_wire2(4, 61)    <= sub_wire1(61);
	sub_wire2(4, 62)    <= sub_wire1(62);
	sub_wire2(4, 63)    <= sub_wire1(63);
	sub_wire2(4, 64)    <= sub_wire1(64);
	sub_wire2(4, 65)    <= sub_wire1(65);
	sub_wire2(4, 66)    <= sub_wire1(66);
	sub_wire2(4, 67)    <= sub_wire1(67);
	sub_wire2(4, 68)    <= sub_wire1(68);
	sub_wire2(4, 69)    <= sub_wire1(69);
	sub_wire2(4, 70)    <= sub_wire1(70);
	sub_wire2(4, 71)    <= sub_wire1(71);
	sub_wire2(4, 72)    <= sub_wire1(72);
	sub_wire2(4, 73)    <= sub_wire1(73);
	sub_wire2(4, 74)    <= sub_wire1(74);
	sub_wire2(4, 75)    <= sub_wire1(75);
	sub_wire2(4, 76)    <= sub_wire1(76);
	sub_wire2(4, 77)    <= sub_wire1(77);
	sub_wire2(4, 78)    <= sub_wire1(78);
	sub_wire2(4, 79)    <= sub_wire1(79);
	sub_wire2(4, 80)    <= sub_wire1(80);
	sub_wire2(4, 81)    <= sub_wire1(81);
	sub_wire2(4, 82)    <= sub_wire1(82);
	sub_wire2(4, 83)    <= sub_wire1(83);
	sub_wire2(4, 84)    <= sub_wire1(84);
	sub_wire2(4, 85)    <= sub_wire1(85);
	sub_wire2(4, 86)    <= sub_wire1(86);
	sub_wire2(4, 87)    <= sub_wire1(87);
	sub_wire2(4, 88)    <= sub_wire1(88);
	sub_wire2(4, 89)    <= sub_wire1(89);
	sub_wire2(4, 90)    <= sub_wire1(90);
	sub_wire2(4, 91)    <= sub_wire1(91);
	sub_wire2(4, 92)    <= sub_wire1(92);
	sub_wire2(4, 93)    <= sub_wire1(93);
	sub_wire2(4, 94)    <= sub_wire1(94);
	sub_wire2(4, 95)    <= sub_wire1(95);
	sub_wire2(4, 96)    <= sub_wire1(96);
	sub_wire2(4, 97)    <= sub_wire1(97);
	sub_wire2(4, 98)    <= sub_wire1(98);
	sub_wire2(4, 99)    <= sub_wire1(99);
	sub_wire2(4, 100)    <= sub_wire1(100);
	sub_wire2(4, 101)    <= sub_wire1(101);
	sub_wire2(4, 102)    <= sub_wire1(102);
	sub_wire2(4, 103)    <= sub_wire1(103);
	sub_wire2(4, 104)    <= sub_wire1(104);
	sub_wire2(4, 105)    <= sub_wire1(105);
	sub_wire2(4, 106)    <= sub_wire1(106);
	sub_wire2(4, 107)    <= sub_wire1(107);
	sub_wire2(4, 108)    <= sub_wire1(108);
	sub_wire2(4, 109)    <= sub_wire1(109);
	sub_wire2(4, 110)    <= sub_wire1(110);
	sub_wire2(4, 111)    <= sub_wire1(111);
	sub_wire2(4, 112)    <= sub_wire1(112);
	sub_wire2(4, 113)    <= sub_wire1(113);
	sub_wire2(4, 114)    <= sub_wire1(114);
	sub_wire2(4, 115)    <= sub_wire1(115);
	sub_wire2(4, 116)    <= sub_wire1(116);
	sub_wire2(4, 117)    <= sub_wire1(117);
	sub_wire2(4, 118)    <= sub_wire1(118);
	sub_wire2(4, 119)    <= sub_wire1(119);
	sub_wire2(4, 120)    <= sub_wire1(120);
	sub_wire2(4, 121)    <= sub_wire1(121);
	sub_wire2(4, 122)    <= sub_wire1(122);
	sub_wire2(4, 123)    <= sub_wire1(123);
	sub_wire2(4, 124)    <= sub_wire1(124);
	sub_wire2(4, 125)    <= sub_wire1(125);
	sub_wire2(4, 126)    <= sub_wire1(126);
	sub_wire2(4, 127)    <= sub_wire1(127);
	sub_wire2(4, 128)    <= sub_wire1(128);
	sub_wire2(4, 129)    <= sub_wire1(129);
	sub_wire2(4, 130)    <= sub_wire1(130);
	sub_wire2(4, 131)    <= sub_wire1(131);
	sub_wire2(4, 132)    <= sub_wire1(132);
	sub_wire2(4, 133)    <= sub_wire1(133);
	sub_wire2(4, 134)    <= sub_wire1(134);
	sub_wire2(4, 135)    <= sub_wire1(135);
	sub_wire2(4, 136)    <= sub_wire1(136);
	sub_wire2(4, 137)    <= sub_wire1(137);
	sub_wire2(4, 138)    <= sub_wire1(138);
	sub_wire2(4, 139)    <= sub_wire1(139);
	sub_wire2(4, 140)    <= sub_wire1(140);
	sub_wire2(4, 141)    <= sub_wire1(141);
	sub_wire2(4, 142)    <= sub_wire1(142);
	sub_wire2(4, 143)    <= sub_wire1(143);
	sub_wire2(4, 144)    <= sub_wire1(144);
	sub_wire2(4, 145)    <= sub_wire1(145);
	sub_wire2(4, 146)    <= sub_wire1(146);
	sub_wire2(4, 147)    <= sub_wire1(147);
	sub_wire2(4, 148)    <= sub_wire1(148);
	sub_wire2(4, 149)    <= sub_wire1(149);
	sub_wire2(4, 150)    <= sub_wire1(150);
	sub_wire2(4, 151)    <= sub_wire1(151);
	sub_wire2(4, 152)    <= sub_wire1(152);
	sub_wire2(4, 153)    <= sub_wire1(153);
	sub_wire2(4, 154)    <= sub_wire1(154);
	sub_wire2(4, 155)    <= sub_wire1(155);
	sub_wire2(4, 156)    <= sub_wire1(156);
	sub_wire2(4, 157)    <= sub_wire1(157);
	sub_wire2(4, 158)    <= sub_wire1(158);
	sub_wire2(4, 159)    <= sub_wire1(159);
	sub_wire2(4, 160)    <= sub_wire1(160);
	sub_wire2(4, 161)    <= sub_wire1(161);
	sub_wire2(4, 162)    <= sub_wire1(162);
	sub_wire2(4, 163)    <= sub_wire1(163);
	sub_wire2(4, 164)    <= sub_wire1(164);
	sub_wire2(4, 165)    <= sub_wire1(165);
	sub_wire2(4, 166)    <= sub_wire1(166);
	sub_wire2(4, 167)    <= sub_wire1(167);
	sub_wire2(4, 168)    <= sub_wire1(168);
	sub_wire2(4, 169)    <= sub_wire1(169);
	sub_wire2(4, 170)    <= sub_wire1(170);
	sub_wire2(4, 171)    <= sub_wire1(171);
	sub_wire2(4, 172)    <= sub_wire1(172);
	sub_wire2(4, 173)    <= sub_wire1(173);
	sub_wire2(4, 174)    <= sub_wire1(174);
	sub_wire2(4, 175)    <= sub_wire1(175);
	sub_wire2(4, 176)    <= sub_wire1(176);
	sub_wire2(4, 177)    <= sub_wire1(177);
	sub_wire2(4, 178)    <= sub_wire1(178);
	sub_wire2(4, 179)    <= sub_wire1(179);
	sub_wire2(3, 0)    <= sub_wire3(0);
	sub_wire2(3, 1)    <= sub_wire3(1);
	sub_wire2(3, 2)    <= sub_wire3(2);
	sub_wire2(3, 3)    <= sub_wire3(3);
	sub_wire2(3, 4)    <= sub_wire3(4);
	sub_wire2(3, 5)    <= sub_wire3(5);
	sub_wire2(3, 6)    <= sub_wire3(6);
	sub_wire2(3, 7)    <= sub_wire3(7);
	sub_wire2(3, 8)    <= sub_wire3(8);
	sub_wire2(3, 9)    <= sub_wire3(9);
	sub_wire2(3, 10)    <= sub_wire3(10);
	sub_wire2(3, 11)    <= sub_wire3(11);
	sub_wire2(3, 12)    <= sub_wire3(12);
	sub_wire2(3, 13)    <= sub_wire3(13);
	sub_wire2(3, 14)    <= sub_wire3(14);
	sub_wire2(3, 15)    <= sub_wire3(15);
	sub_wire2(3, 16)    <= sub_wire3(16);
	sub_wire2(3, 17)    <= sub_wire3(17);
	sub_wire2(3, 18)    <= sub_wire3(18);
	sub_wire2(3, 19)    <= sub_wire3(19);
	sub_wire2(3, 20)    <= sub_wire3(20);
	sub_wire2(3, 21)    <= sub_wire3(21);
	sub_wire2(3, 22)    <= sub_wire3(22);
	sub_wire2(3, 23)    <= sub_wire3(23);
	sub_wire2(3, 24)    <= sub_wire3(24);
	sub_wire2(3, 25)    <= sub_wire3(25);
	sub_wire2(3, 26)    <= sub_wire3(26);
	sub_wire2(3, 27)    <= sub_wire3(27);
	sub_wire2(3, 28)    <= sub_wire3(28);
	sub_wire2(3, 29)    <= sub_wire3(29);
	sub_wire2(3, 30)    <= sub_wire3(30);
	sub_wire2(3, 31)    <= sub_wire3(31);
	sub_wire2(3, 32)    <= sub_wire3(32);
	sub_wire2(3, 33)    <= sub_wire3(33);
	sub_wire2(3, 34)    <= sub_wire3(34);
	sub_wire2(3, 35)    <= sub_wire3(35);
	sub_wire2(3, 36)    <= sub_wire3(36);
	sub_wire2(3, 37)    <= sub_wire3(37);
	sub_wire2(3, 38)    <= sub_wire3(38);
	sub_wire2(3, 39)    <= sub_wire3(39);
	sub_wire2(3, 40)    <= sub_wire3(40);
	sub_wire2(3, 41)    <= sub_wire3(41);
	sub_wire2(3, 42)    <= sub_wire3(42);
	sub_wire2(3, 43)    <= sub_wire3(43);
	sub_wire2(3, 44)    <= sub_wire3(44);
	sub_wire2(3, 45)    <= sub_wire3(45);
	sub_wire2(3, 46)    <= sub_wire3(46);
	sub_wire2(3, 47)    <= sub_wire3(47);
	sub_wire2(3, 48)    <= sub_wire3(48);
	sub_wire2(3, 49)    <= sub_wire3(49);
	sub_wire2(3, 50)    <= sub_wire3(50);
	sub_wire2(3, 51)    <= sub_wire3(51);
	sub_wire2(3, 52)    <= sub_wire3(52);
	sub_wire2(3, 53)    <= sub_wire3(53);
	sub_wire2(3, 54)    <= sub_wire3(54);
	sub_wire2(3, 55)    <= sub_wire3(55);
	sub_wire2(3, 56)    <= sub_wire3(56);
	sub_wire2(3, 57)    <= sub_wire3(57);
	sub_wire2(3, 58)    <= sub_wire3(58);
	sub_wire2(3, 59)    <= sub_wire3(59);
	sub_wire2(3, 60)    <= sub_wire3(60);
	sub_wire2(3, 61)    <= sub_wire3(61);
	sub_wire2(3, 62)    <= sub_wire3(62);
	sub_wire2(3, 63)    <= sub_wire3(63);
	sub_wire2(3, 64)    <= sub_wire3(64);
	sub_wire2(3, 65)    <= sub_wire3(65);
	sub_wire2(3, 66)    <= sub_wire3(66);
	sub_wire2(3, 67)    <= sub_wire3(67);
	sub_wire2(3, 68)    <= sub_wire3(68);
	sub_wire2(3, 69)    <= sub_wire3(69);
	sub_wire2(3, 70)    <= sub_wire3(70);
	sub_wire2(3, 71)    <= sub_wire3(71);
	sub_wire2(3, 72)    <= sub_wire3(72);
	sub_wire2(3, 73)    <= sub_wire3(73);
	sub_wire2(3, 74)    <= sub_wire3(74);
	sub_wire2(3, 75)    <= sub_wire3(75);
	sub_wire2(3, 76)    <= sub_wire3(76);
	sub_wire2(3, 77)    <= sub_wire3(77);
	sub_wire2(3, 78)    <= sub_wire3(78);
	sub_wire2(3, 79)    <= sub_wire3(79);
	sub_wire2(3, 80)    <= sub_wire3(80);
	sub_wire2(3, 81)    <= sub_wire3(81);
	sub_wire2(3, 82)    <= sub_wire3(82);
	sub_wire2(3, 83)    <= sub_wire3(83);
	sub_wire2(3, 84)    <= sub_wire3(84);
	sub_wire2(3, 85)    <= sub_wire3(85);
	sub_wire2(3, 86)    <= sub_wire3(86);
	sub_wire2(3, 87)    <= sub_wire3(87);
	sub_wire2(3, 88)    <= sub_wire3(88);
	sub_wire2(3, 89)    <= sub_wire3(89);
	sub_wire2(3, 90)    <= sub_wire3(90);
	sub_wire2(3, 91)    <= sub_wire3(91);
	sub_wire2(3, 92)    <= sub_wire3(92);
	sub_wire2(3, 93)    <= sub_wire3(93);
	sub_wire2(3, 94)    <= sub_wire3(94);
	sub_wire2(3, 95)    <= sub_wire3(95);
	sub_wire2(3, 96)    <= sub_wire3(96);
	sub_wire2(3, 97)    <= sub_wire3(97);
	sub_wire2(3, 98)    <= sub_wire3(98);
	sub_wire2(3, 99)    <= sub_wire3(99);
	sub_wire2(3, 100)    <= sub_wire3(100);
	sub_wire2(3, 101)    <= sub_wire3(101);
	sub_wire2(3, 102)    <= sub_wire3(102);
	sub_wire2(3, 103)    <= sub_wire3(103);
	sub_wire2(3, 104)    <= sub_wire3(104);
	sub_wire2(3, 105)    <= sub_wire3(105);
	sub_wire2(3, 106)    <= sub_wire3(106);
	sub_wire2(3, 107)    <= sub_wire3(107);
	sub_wire2(3, 108)    <= sub_wire3(108);
	sub_wire2(3, 109)    <= sub_wire3(109);
	sub_wire2(3, 110)    <= sub_wire3(110);
	sub_wire2(3, 111)    <= sub_wire3(111);
	sub_wire2(3, 112)    <= sub_wire3(112);
	sub_wire2(3, 113)    <= sub_wire3(113);
	sub_wire2(3, 114)    <= sub_wire3(114);
	sub_wire2(3, 115)    <= sub_wire3(115);
	sub_wire2(3, 116)    <= sub_wire3(116);
	sub_wire2(3, 117)    <= sub_wire3(117);
	sub_wire2(3, 118)    <= sub_wire3(118);
	sub_wire2(3, 119)    <= sub_wire3(119);
	sub_wire2(3, 120)    <= sub_wire3(120);
	sub_wire2(3, 121)    <= sub_wire3(121);
	sub_wire2(3, 122)    <= sub_wire3(122);
	sub_wire2(3, 123)    <= sub_wire3(123);
	sub_wire2(3, 124)    <= sub_wire3(124);
	sub_wire2(3, 125)    <= sub_wire3(125);
	sub_wire2(3, 126)    <= sub_wire3(126);
	sub_wire2(3, 127)    <= sub_wire3(127);
	sub_wire2(3, 128)    <= sub_wire3(128);
	sub_wire2(3, 129)    <= sub_wire3(129);
	sub_wire2(3, 130)    <= sub_wire3(130);
	sub_wire2(3, 131)    <= sub_wire3(131);
	sub_wire2(3, 132)    <= sub_wire3(132);
	sub_wire2(3, 133)    <= sub_wire3(133);
	sub_wire2(3, 134)    <= sub_wire3(134);
	sub_wire2(3, 135)    <= sub_wire3(135);
	sub_wire2(3, 136)    <= sub_wire3(136);
	sub_wire2(3, 137)    <= sub_wire3(137);
	sub_wire2(3, 138)    <= sub_wire3(138);
	sub_wire2(3, 139)    <= sub_wire3(139);
	sub_wire2(3, 140)    <= sub_wire3(140);
	sub_wire2(3, 141)    <= sub_wire3(141);
	sub_wire2(3, 142)    <= sub_wire3(142);
	sub_wire2(3, 143)    <= sub_wire3(143);
	sub_wire2(3, 144)    <= sub_wire3(144);
	sub_wire2(3, 145)    <= sub_wire3(145);
	sub_wire2(3, 146)    <= sub_wire3(146);
	sub_wire2(3, 147)    <= sub_wire3(147);
	sub_wire2(3, 148)    <= sub_wire3(148);
	sub_wire2(3, 149)    <= sub_wire3(149);
	sub_wire2(3, 150)    <= sub_wire3(150);
	sub_wire2(3, 151)    <= sub_wire3(151);
	sub_wire2(3, 152)    <= sub_wire3(152);
	sub_wire2(3, 153)    <= sub_wire3(153);
	sub_wire2(3, 154)    <= sub_wire3(154);
	sub_wire2(3, 155)    <= sub_wire3(155);
	sub_wire2(3, 156)    <= sub_wire3(156);
	sub_wire2(3, 157)    <= sub_wire3(157);
	sub_wire2(3, 158)    <= sub_wire3(158);
	sub_wire2(3, 159)    <= sub_wire3(159);
	sub_wire2(3, 160)    <= sub_wire3(160);
	sub_wire2(3, 161)    <= sub_wire3(161);
	sub_wire2(3, 162)    <= sub_wire3(162);
	sub_wire2(3, 163)    <= sub_wire3(163);
	sub_wire2(3, 164)    <= sub_wire3(164);
	sub_wire2(3, 165)    <= sub_wire3(165);
	sub_wire2(3, 166)    <= sub_wire3(166);
	sub_wire2(3, 167)    <= sub_wire3(167);
	sub_wire2(3, 168)    <= sub_wire3(168);
	sub_wire2(3, 169)    <= sub_wire3(169);
	sub_wire2(3, 170)    <= sub_wire3(170);
	sub_wire2(3, 171)    <= sub_wire3(171);
	sub_wire2(3, 172)    <= sub_wire3(172);
	sub_wire2(3, 173)    <= sub_wire3(173);
	sub_wire2(3, 174)    <= sub_wire3(174);
	sub_wire2(3, 175)    <= sub_wire3(175);
	sub_wire2(3, 176)    <= sub_wire3(176);
	sub_wire2(3, 177)    <= sub_wire3(177);
	sub_wire2(3, 178)    <= sub_wire3(178);
	sub_wire2(3, 179)    <= sub_wire3(179);
	sub_wire2(2, 0)    <= sub_wire4(0);
	sub_wire2(2, 1)    <= sub_wire4(1);
	sub_wire2(2, 2)    <= sub_wire4(2);
	sub_wire2(2, 3)    <= sub_wire4(3);
	sub_wire2(2, 4)    <= sub_wire4(4);
	sub_wire2(2, 5)    <= sub_wire4(5);
	sub_wire2(2, 6)    <= sub_wire4(6);
	sub_wire2(2, 7)    <= sub_wire4(7);
	sub_wire2(2, 8)    <= sub_wire4(8);
	sub_wire2(2, 9)    <= sub_wire4(9);
	sub_wire2(2, 10)    <= sub_wire4(10);
	sub_wire2(2, 11)    <= sub_wire4(11);
	sub_wire2(2, 12)    <= sub_wire4(12);
	sub_wire2(2, 13)    <= sub_wire4(13);
	sub_wire2(2, 14)    <= sub_wire4(14);
	sub_wire2(2, 15)    <= sub_wire4(15);
	sub_wire2(2, 16)    <= sub_wire4(16);
	sub_wire2(2, 17)    <= sub_wire4(17);
	sub_wire2(2, 18)    <= sub_wire4(18);
	sub_wire2(2, 19)    <= sub_wire4(19);
	sub_wire2(2, 20)    <= sub_wire4(20);
	sub_wire2(2, 21)    <= sub_wire4(21);
	sub_wire2(2, 22)    <= sub_wire4(22);
	sub_wire2(2, 23)    <= sub_wire4(23);
	sub_wire2(2, 24)    <= sub_wire4(24);
	sub_wire2(2, 25)    <= sub_wire4(25);
	sub_wire2(2, 26)    <= sub_wire4(26);
	sub_wire2(2, 27)    <= sub_wire4(27);
	sub_wire2(2, 28)    <= sub_wire4(28);
	sub_wire2(2, 29)    <= sub_wire4(29);
	sub_wire2(2, 30)    <= sub_wire4(30);
	sub_wire2(2, 31)    <= sub_wire4(31);
	sub_wire2(2, 32)    <= sub_wire4(32);
	sub_wire2(2, 33)    <= sub_wire4(33);
	sub_wire2(2, 34)    <= sub_wire4(34);
	sub_wire2(2, 35)    <= sub_wire4(35);
	sub_wire2(2, 36)    <= sub_wire4(36);
	sub_wire2(2, 37)    <= sub_wire4(37);
	sub_wire2(2, 38)    <= sub_wire4(38);
	sub_wire2(2, 39)    <= sub_wire4(39);
	sub_wire2(2, 40)    <= sub_wire4(40);
	sub_wire2(2, 41)    <= sub_wire4(41);
	sub_wire2(2, 42)    <= sub_wire4(42);
	sub_wire2(2, 43)    <= sub_wire4(43);
	sub_wire2(2, 44)    <= sub_wire4(44);
	sub_wire2(2, 45)    <= sub_wire4(45);
	sub_wire2(2, 46)    <= sub_wire4(46);
	sub_wire2(2, 47)    <= sub_wire4(47);
	sub_wire2(2, 48)    <= sub_wire4(48);
	sub_wire2(2, 49)    <= sub_wire4(49);
	sub_wire2(2, 50)    <= sub_wire4(50);
	sub_wire2(2, 51)    <= sub_wire4(51);
	sub_wire2(2, 52)    <= sub_wire4(52);
	sub_wire2(2, 53)    <= sub_wire4(53);
	sub_wire2(2, 54)    <= sub_wire4(54);
	sub_wire2(2, 55)    <= sub_wire4(55);
	sub_wire2(2, 56)    <= sub_wire4(56);
	sub_wire2(2, 57)    <= sub_wire4(57);
	sub_wire2(2, 58)    <= sub_wire4(58);
	sub_wire2(2, 59)    <= sub_wire4(59);
	sub_wire2(2, 60)    <= sub_wire4(60);
	sub_wire2(2, 61)    <= sub_wire4(61);
	sub_wire2(2, 62)    <= sub_wire4(62);
	sub_wire2(2, 63)    <= sub_wire4(63);
	sub_wire2(2, 64)    <= sub_wire4(64);
	sub_wire2(2, 65)    <= sub_wire4(65);
	sub_wire2(2, 66)    <= sub_wire4(66);
	sub_wire2(2, 67)    <= sub_wire4(67);
	sub_wire2(2, 68)    <= sub_wire4(68);
	sub_wire2(2, 69)    <= sub_wire4(69);
	sub_wire2(2, 70)    <= sub_wire4(70);
	sub_wire2(2, 71)    <= sub_wire4(71);
	sub_wire2(2, 72)    <= sub_wire4(72);
	sub_wire2(2, 73)    <= sub_wire4(73);
	sub_wire2(2, 74)    <= sub_wire4(74);
	sub_wire2(2, 75)    <= sub_wire4(75);
	sub_wire2(2, 76)    <= sub_wire4(76);
	sub_wire2(2, 77)    <= sub_wire4(77);
	sub_wire2(2, 78)    <= sub_wire4(78);
	sub_wire2(2, 79)    <= sub_wire4(79);
	sub_wire2(2, 80)    <= sub_wire4(80);
	sub_wire2(2, 81)    <= sub_wire4(81);
	sub_wire2(2, 82)    <= sub_wire4(82);
	sub_wire2(2, 83)    <= sub_wire4(83);
	sub_wire2(2, 84)    <= sub_wire4(84);
	sub_wire2(2, 85)    <= sub_wire4(85);
	sub_wire2(2, 86)    <= sub_wire4(86);
	sub_wire2(2, 87)    <= sub_wire4(87);
	sub_wire2(2, 88)    <= sub_wire4(88);
	sub_wire2(2, 89)    <= sub_wire4(89);
	sub_wire2(2, 90)    <= sub_wire4(90);
	sub_wire2(2, 91)    <= sub_wire4(91);
	sub_wire2(2, 92)    <= sub_wire4(92);
	sub_wire2(2, 93)    <= sub_wire4(93);
	sub_wire2(2, 94)    <= sub_wire4(94);
	sub_wire2(2, 95)    <= sub_wire4(95);
	sub_wire2(2, 96)    <= sub_wire4(96);
	sub_wire2(2, 97)    <= sub_wire4(97);
	sub_wire2(2, 98)    <= sub_wire4(98);
	sub_wire2(2, 99)    <= sub_wire4(99);
	sub_wire2(2, 100)    <= sub_wire4(100);
	sub_wire2(2, 101)    <= sub_wire4(101);
	sub_wire2(2, 102)    <= sub_wire4(102);
	sub_wire2(2, 103)    <= sub_wire4(103);
	sub_wire2(2, 104)    <= sub_wire4(104);
	sub_wire2(2, 105)    <= sub_wire4(105);
	sub_wire2(2, 106)    <= sub_wire4(106);
	sub_wire2(2, 107)    <= sub_wire4(107);
	sub_wire2(2, 108)    <= sub_wire4(108);
	sub_wire2(2, 109)    <= sub_wire4(109);
	sub_wire2(2, 110)    <= sub_wire4(110);
	sub_wire2(2, 111)    <= sub_wire4(111);
	sub_wire2(2, 112)    <= sub_wire4(112);
	sub_wire2(2, 113)    <= sub_wire4(113);
	sub_wire2(2, 114)    <= sub_wire4(114);
	sub_wire2(2, 115)    <= sub_wire4(115);
	sub_wire2(2, 116)    <= sub_wire4(116);
	sub_wire2(2, 117)    <= sub_wire4(117);
	sub_wire2(2, 118)    <= sub_wire4(118);
	sub_wire2(2, 119)    <= sub_wire4(119);
	sub_wire2(2, 120)    <= sub_wire4(120);
	sub_wire2(2, 121)    <= sub_wire4(121);
	sub_wire2(2, 122)    <= sub_wire4(122);
	sub_wire2(2, 123)    <= sub_wire4(123);
	sub_wire2(2, 124)    <= sub_wire4(124);
	sub_wire2(2, 125)    <= sub_wire4(125);
	sub_wire2(2, 126)    <= sub_wire4(126);
	sub_wire2(2, 127)    <= sub_wire4(127);
	sub_wire2(2, 128)    <= sub_wire4(128);
	sub_wire2(2, 129)    <= sub_wire4(129);
	sub_wire2(2, 130)    <= sub_wire4(130);
	sub_wire2(2, 131)    <= sub_wire4(131);
	sub_wire2(2, 132)    <= sub_wire4(132);
	sub_wire2(2, 133)    <= sub_wire4(133);
	sub_wire2(2, 134)    <= sub_wire4(134);
	sub_wire2(2, 135)    <= sub_wire4(135);
	sub_wire2(2, 136)    <= sub_wire4(136);
	sub_wire2(2, 137)    <= sub_wire4(137);
	sub_wire2(2, 138)    <= sub_wire4(138);
	sub_wire2(2, 139)    <= sub_wire4(139);
	sub_wire2(2, 140)    <= sub_wire4(140);
	sub_wire2(2, 141)    <= sub_wire4(141);
	sub_wire2(2, 142)    <= sub_wire4(142);
	sub_wire2(2, 143)    <= sub_wire4(143);
	sub_wire2(2, 144)    <= sub_wire4(144);
	sub_wire2(2, 145)    <= sub_wire4(145);
	sub_wire2(2, 146)    <= sub_wire4(146);
	sub_wire2(2, 147)    <= sub_wire4(147);
	sub_wire2(2, 148)    <= sub_wire4(148);
	sub_wire2(2, 149)    <= sub_wire4(149);
	sub_wire2(2, 150)    <= sub_wire4(150);
	sub_wire2(2, 151)    <= sub_wire4(151);
	sub_wire2(2, 152)    <= sub_wire4(152);
	sub_wire2(2, 153)    <= sub_wire4(153);
	sub_wire2(2, 154)    <= sub_wire4(154);
	sub_wire2(2, 155)    <= sub_wire4(155);
	sub_wire2(2, 156)    <= sub_wire4(156);
	sub_wire2(2, 157)    <= sub_wire4(157);
	sub_wire2(2, 158)    <= sub_wire4(158);
	sub_wire2(2, 159)    <= sub_wire4(159);
	sub_wire2(2, 160)    <= sub_wire4(160);
	sub_wire2(2, 161)    <= sub_wire4(161);
	sub_wire2(2, 162)    <= sub_wire4(162);
	sub_wire2(2, 163)    <= sub_wire4(163);
	sub_wire2(2, 164)    <= sub_wire4(164);
	sub_wire2(2, 165)    <= sub_wire4(165);
	sub_wire2(2, 166)    <= sub_wire4(166);
	sub_wire2(2, 167)    <= sub_wire4(167);
	sub_wire2(2, 168)    <= sub_wire4(168);
	sub_wire2(2, 169)    <= sub_wire4(169);
	sub_wire2(2, 170)    <= sub_wire4(170);
	sub_wire2(2, 171)    <= sub_wire4(171);
	sub_wire2(2, 172)    <= sub_wire4(172);
	sub_wire2(2, 173)    <= sub_wire4(173);
	sub_wire2(2, 174)    <= sub_wire4(174);
	sub_wire2(2, 175)    <= sub_wire4(175);
	sub_wire2(2, 176)    <= sub_wire4(176);
	sub_wire2(2, 177)    <= sub_wire4(177);
	sub_wire2(2, 178)    <= sub_wire4(178);
	sub_wire2(2, 179)    <= sub_wire4(179);
	sub_wire2(1, 0)    <= sub_wire5(0);
	sub_wire2(1, 1)    <= sub_wire5(1);
	sub_wire2(1, 2)    <= sub_wire5(2);
	sub_wire2(1, 3)    <= sub_wire5(3);
	sub_wire2(1, 4)    <= sub_wire5(4);
	sub_wire2(1, 5)    <= sub_wire5(5);
	sub_wire2(1, 6)    <= sub_wire5(6);
	sub_wire2(1, 7)    <= sub_wire5(7);
	sub_wire2(1, 8)    <= sub_wire5(8);
	sub_wire2(1, 9)    <= sub_wire5(9);
	sub_wire2(1, 10)    <= sub_wire5(10);
	sub_wire2(1, 11)    <= sub_wire5(11);
	sub_wire2(1, 12)    <= sub_wire5(12);
	sub_wire2(1, 13)    <= sub_wire5(13);
	sub_wire2(1, 14)    <= sub_wire5(14);
	sub_wire2(1, 15)    <= sub_wire5(15);
	sub_wire2(1, 16)    <= sub_wire5(16);
	sub_wire2(1, 17)    <= sub_wire5(17);
	sub_wire2(1, 18)    <= sub_wire5(18);
	sub_wire2(1, 19)    <= sub_wire5(19);
	sub_wire2(1, 20)    <= sub_wire5(20);
	sub_wire2(1, 21)    <= sub_wire5(21);
	sub_wire2(1, 22)    <= sub_wire5(22);
	sub_wire2(1, 23)    <= sub_wire5(23);
	sub_wire2(1, 24)    <= sub_wire5(24);
	sub_wire2(1, 25)    <= sub_wire5(25);
	sub_wire2(1, 26)    <= sub_wire5(26);
	sub_wire2(1, 27)    <= sub_wire5(27);
	sub_wire2(1, 28)    <= sub_wire5(28);
	sub_wire2(1, 29)    <= sub_wire5(29);
	sub_wire2(1, 30)    <= sub_wire5(30);
	sub_wire2(1, 31)    <= sub_wire5(31);
	sub_wire2(1, 32)    <= sub_wire5(32);
	sub_wire2(1, 33)    <= sub_wire5(33);
	sub_wire2(1, 34)    <= sub_wire5(34);
	sub_wire2(1, 35)    <= sub_wire5(35);
	sub_wire2(1, 36)    <= sub_wire5(36);
	sub_wire2(1, 37)    <= sub_wire5(37);
	sub_wire2(1, 38)    <= sub_wire5(38);
	sub_wire2(1, 39)    <= sub_wire5(39);
	sub_wire2(1, 40)    <= sub_wire5(40);
	sub_wire2(1, 41)    <= sub_wire5(41);
	sub_wire2(1, 42)    <= sub_wire5(42);
	sub_wire2(1, 43)    <= sub_wire5(43);
	sub_wire2(1, 44)    <= sub_wire5(44);
	sub_wire2(1, 45)    <= sub_wire5(45);
	sub_wire2(1, 46)    <= sub_wire5(46);
	sub_wire2(1, 47)    <= sub_wire5(47);
	sub_wire2(1, 48)    <= sub_wire5(48);
	sub_wire2(1, 49)    <= sub_wire5(49);
	sub_wire2(1, 50)    <= sub_wire5(50);
	sub_wire2(1, 51)    <= sub_wire5(51);
	sub_wire2(1, 52)    <= sub_wire5(52);
	sub_wire2(1, 53)    <= sub_wire5(53);
	sub_wire2(1, 54)    <= sub_wire5(54);
	sub_wire2(1, 55)    <= sub_wire5(55);
	sub_wire2(1, 56)    <= sub_wire5(56);
	sub_wire2(1, 57)    <= sub_wire5(57);
	sub_wire2(1, 58)    <= sub_wire5(58);
	sub_wire2(1, 59)    <= sub_wire5(59);
	sub_wire2(1, 60)    <= sub_wire5(60);
	sub_wire2(1, 61)    <= sub_wire5(61);
	sub_wire2(1, 62)    <= sub_wire5(62);
	sub_wire2(1, 63)    <= sub_wire5(63);
	sub_wire2(1, 64)    <= sub_wire5(64);
	sub_wire2(1, 65)    <= sub_wire5(65);
	sub_wire2(1, 66)    <= sub_wire5(66);
	sub_wire2(1, 67)    <= sub_wire5(67);
	sub_wire2(1, 68)    <= sub_wire5(68);
	sub_wire2(1, 69)    <= sub_wire5(69);
	sub_wire2(1, 70)    <= sub_wire5(70);
	sub_wire2(1, 71)    <= sub_wire5(71);
	sub_wire2(1, 72)    <= sub_wire5(72);
	sub_wire2(1, 73)    <= sub_wire5(73);
	sub_wire2(1, 74)    <= sub_wire5(74);
	sub_wire2(1, 75)    <= sub_wire5(75);
	sub_wire2(1, 76)    <= sub_wire5(76);
	sub_wire2(1, 77)    <= sub_wire5(77);
	sub_wire2(1, 78)    <= sub_wire5(78);
	sub_wire2(1, 79)    <= sub_wire5(79);
	sub_wire2(1, 80)    <= sub_wire5(80);
	sub_wire2(1, 81)    <= sub_wire5(81);
	sub_wire2(1, 82)    <= sub_wire5(82);
	sub_wire2(1, 83)    <= sub_wire5(83);
	sub_wire2(1, 84)    <= sub_wire5(84);
	sub_wire2(1, 85)    <= sub_wire5(85);
	sub_wire2(1, 86)    <= sub_wire5(86);
	sub_wire2(1, 87)    <= sub_wire5(87);
	sub_wire2(1, 88)    <= sub_wire5(88);
	sub_wire2(1, 89)    <= sub_wire5(89);
	sub_wire2(1, 90)    <= sub_wire5(90);
	sub_wire2(1, 91)    <= sub_wire5(91);
	sub_wire2(1, 92)    <= sub_wire5(92);
	sub_wire2(1, 93)    <= sub_wire5(93);
	sub_wire2(1, 94)    <= sub_wire5(94);
	sub_wire2(1, 95)    <= sub_wire5(95);
	sub_wire2(1, 96)    <= sub_wire5(96);
	sub_wire2(1, 97)    <= sub_wire5(97);
	sub_wire2(1, 98)    <= sub_wire5(98);
	sub_wire2(1, 99)    <= sub_wire5(99);
	sub_wire2(1, 100)    <= sub_wire5(100);
	sub_wire2(1, 101)    <= sub_wire5(101);
	sub_wire2(1, 102)    <= sub_wire5(102);
	sub_wire2(1, 103)    <= sub_wire5(103);
	sub_wire2(1, 104)    <= sub_wire5(104);
	sub_wire2(1, 105)    <= sub_wire5(105);
	sub_wire2(1, 106)    <= sub_wire5(106);
	sub_wire2(1, 107)    <= sub_wire5(107);
	sub_wire2(1, 108)    <= sub_wire5(108);
	sub_wire2(1, 109)    <= sub_wire5(109);
	sub_wire2(1, 110)    <= sub_wire5(110);
	sub_wire2(1, 111)    <= sub_wire5(111);
	sub_wire2(1, 112)    <= sub_wire5(112);
	sub_wire2(1, 113)    <= sub_wire5(113);
	sub_wire2(1, 114)    <= sub_wire5(114);
	sub_wire2(1, 115)    <= sub_wire5(115);
	sub_wire2(1, 116)    <= sub_wire5(116);
	sub_wire2(1, 117)    <= sub_wire5(117);
	sub_wire2(1, 118)    <= sub_wire5(118);
	sub_wire2(1, 119)    <= sub_wire5(119);
	sub_wire2(1, 120)    <= sub_wire5(120);
	sub_wire2(1, 121)    <= sub_wire5(121);
	sub_wire2(1, 122)    <= sub_wire5(122);
	sub_wire2(1, 123)    <= sub_wire5(123);
	sub_wire2(1, 124)    <= sub_wire5(124);
	sub_wire2(1, 125)    <= sub_wire5(125);
	sub_wire2(1, 126)    <= sub_wire5(126);
	sub_wire2(1, 127)    <= sub_wire5(127);
	sub_wire2(1, 128)    <= sub_wire5(128);
	sub_wire2(1, 129)    <= sub_wire5(129);
	sub_wire2(1, 130)    <= sub_wire5(130);
	sub_wire2(1, 131)    <= sub_wire5(131);
	sub_wire2(1, 132)    <= sub_wire5(132);
	sub_wire2(1, 133)    <= sub_wire5(133);
	sub_wire2(1, 134)    <= sub_wire5(134);
	sub_wire2(1, 135)    <= sub_wire5(135);
	sub_wire2(1, 136)    <= sub_wire5(136);
	sub_wire2(1, 137)    <= sub_wire5(137);
	sub_wire2(1, 138)    <= sub_wire5(138);
	sub_wire2(1, 139)    <= sub_wire5(139);
	sub_wire2(1, 140)    <= sub_wire5(140);
	sub_wire2(1, 141)    <= sub_wire5(141);
	sub_wire2(1, 142)    <= sub_wire5(142);
	sub_wire2(1, 143)    <= sub_wire5(143);
	sub_wire2(1, 144)    <= sub_wire5(144);
	sub_wire2(1, 145)    <= sub_wire5(145);
	sub_wire2(1, 146)    <= sub_wire5(146);
	sub_wire2(1, 147)    <= sub_wire5(147);
	sub_wire2(1, 148)    <= sub_wire5(148);
	sub_wire2(1, 149)    <= sub_wire5(149);
	sub_wire2(1, 150)    <= sub_wire5(150);
	sub_wire2(1, 151)    <= sub_wire5(151);
	sub_wire2(1, 152)    <= sub_wire5(152);
	sub_wire2(1, 153)    <= sub_wire5(153);
	sub_wire2(1, 154)    <= sub_wire5(154);
	sub_wire2(1, 155)    <= sub_wire5(155);
	sub_wire2(1, 156)    <= sub_wire5(156);
	sub_wire2(1, 157)    <= sub_wire5(157);
	sub_wire2(1, 158)    <= sub_wire5(158);
	sub_wire2(1, 159)    <= sub_wire5(159);
	sub_wire2(1, 160)    <= sub_wire5(160);
	sub_wire2(1, 161)    <= sub_wire5(161);
	sub_wire2(1, 162)    <= sub_wire5(162);
	sub_wire2(1, 163)    <= sub_wire5(163);
	sub_wire2(1, 164)    <= sub_wire5(164);
	sub_wire2(1, 165)    <= sub_wire5(165);
	sub_wire2(1, 166)    <= sub_wire5(166);
	sub_wire2(1, 167)    <= sub_wire5(167);
	sub_wire2(1, 168)    <= sub_wire5(168);
	sub_wire2(1, 169)    <= sub_wire5(169);
	sub_wire2(1, 170)    <= sub_wire5(170);
	sub_wire2(1, 171)    <= sub_wire5(171);
	sub_wire2(1, 172)    <= sub_wire5(172);
	sub_wire2(1, 173)    <= sub_wire5(173);
	sub_wire2(1, 174)    <= sub_wire5(174);
	sub_wire2(1, 175)    <= sub_wire5(175);
	sub_wire2(1, 176)    <= sub_wire5(176);
	sub_wire2(1, 177)    <= sub_wire5(177);
	sub_wire2(1, 178)    <= sub_wire5(178);
	sub_wire2(1, 179)    <= sub_wire5(179);
	sub_wire2(0, 0)    <= sub_wire6(0);
	sub_wire2(0, 1)    <= sub_wire6(1);
	sub_wire2(0, 2)    <= sub_wire6(2);
	sub_wire2(0, 3)    <= sub_wire6(3);
	sub_wire2(0, 4)    <= sub_wire6(4);
	sub_wire2(0, 5)    <= sub_wire6(5);
	sub_wire2(0, 6)    <= sub_wire6(6);
	sub_wire2(0, 7)    <= sub_wire6(7);
	sub_wire2(0, 8)    <= sub_wire6(8);
	sub_wire2(0, 9)    <= sub_wire6(9);
	sub_wire2(0, 10)    <= sub_wire6(10);
	sub_wire2(0, 11)    <= sub_wire6(11);
	sub_wire2(0, 12)    <= sub_wire6(12);
	sub_wire2(0, 13)    <= sub_wire6(13);
	sub_wire2(0, 14)    <= sub_wire6(14);
	sub_wire2(0, 15)    <= sub_wire6(15);
	sub_wire2(0, 16)    <= sub_wire6(16);
	sub_wire2(0, 17)    <= sub_wire6(17);
	sub_wire2(0, 18)    <= sub_wire6(18);
	sub_wire2(0, 19)    <= sub_wire6(19);
	sub_wire2(0, 20)    <= sub_wire6(20);
	sub_wire2(0, 21)    <= sub_wire6(21);
	sub_wire2(0, 22)    <= sub_wire6(22);
	sub_wire2(0, 23)    <= sub_wire6(23);
	sub_wire2(0, 24)    <= sub_wire6(24);
	sub_wire2(0, 25)    <= sub_wire6(25);
	sub_wire2(0, 26)    <= sub_wire6(26);
	sub_wire2(0, 27)    <= sub_wire6(27);
	sub_wire2(0, 28)    <= sub_wire6(28);
	sub_wire2(0, 29)    <= sub_wire6(29);
	sub_wire2(0, 30)    <= sub_wire6(30);
	sub_wire2(0, 31)    <= sub_wire6(31);
	sub_wire2(0, 32)    <= sub_wire6(32);
	sub_wire2(0, 33)    <= sub_wire6(33);
	sub_wire2(0, 34)    <= sub_wire6(34);
	sub_wire2(0, 35)    <= sub_wire6(35);
	sub_wire2(0, 36)    <= sub_wire6(36);
	sub_wire2(0, 37)    <= sub_wire6(37);
	sub_wire2(0, 38)    <= sub_wire6(38);
	sub_wire2(0, 39)    <= sub_wire6(39);
	sub_wire2(0, 40)    <= sub_wire6(40);
	sub_wire2(0, 41)    <= sub_wire6(41);
	sub_wire2(0, 42)    <= sub_wire6(42);
	sub_wire2(0, 43)    <= sub_wire6(43);
	sub_wire2(0, 44)    <= sub_wire6(44);
	sub_wire2(0, 45)    <= sub_wire6(45);
	sub_wire2(0, 46)    <= sub_wire6(46);
	sub_wire2(0, 47)    <= sub_wire6(47);
	sub_wire2(0, 48)    <= sub_wire6(48);
	sub_wire2(0, 49)    <= sub_wire6(49);
	sub_wire2(0, 50)    <= sub_wire6(50);
	sub_wire2(0, 51)    <= sub_wire6(51);
	sub_wire2(0, 52)    <= sub_wire6(52);
	sub_wire2(0, 53)    <= sub_wire6(53);
	sub_wire2(0, 54)    <= sub_wire6(54);
	sub_wire2(0, 55)    <= sub_wire6(55);
	sub_wire2(0, 56)    <= sub_wire6(56);
	sub_wire2(0, 57)    <= sub_wire6(57);
	sub_wire2(0, 58)    <= sub_wire6(58);
	sub_wire2(0, 59)    <= sub_wire6(59);
	sub_wire2(0, 60)    <= sub_wire6(60);
	sub_wire2(0, 61)    <= sub_wire6(61);
	sub_wire2(0, 62)    <= sub_wire6(62);
	sub_wire2(0, 63)    <= sub_wire6(63);
	sub_wire2(0, 64)    <= sub_wire6(64);
	sub_wire2(0, 65)    <= sub_wire6(65);
	sub_wire2(0, 66)    <= sub_wire6(66);
	sub_wire2(0, 67)    <= sub_wire6(67);
	sub_wire2(0, 68)    <= sub_wire6(68);
	sub_wire2(0, 69)    <= sub_wire6(69);
	sub_wire2(0, 70)    <= sub_wire6(70);
	sub_wire2(0, 71)    <= sub_wire6(71);
	sub_wire2(0, 72)    <= sub_wire6(72);
	sub_wire2(0, 73)    <= sub_wire6(73);
	sub_wire2(0, 74)    <= sub_wire6(74);
	sub_wire2(0, 75)    <= sub_wire6(75);
	sub_wire2(0, 76)    <= sub_wire6(76);
	sub_wire2(0, 77)    <= sub_wire6(77);
	sub_wire2(0, 78)    <= sub_wire6(78);
	sub_wire2(0, 79)    <= sub_wire6(79);
	sub_wire2(0, 80)    <= sub_wire6(80);
	sub_wire2(0, 81)    <= sub_wire6(81);
	sub_wire2(0, 82)    <= sub_wire6(82);
	sub_wire2(0, 83)    <= sub_wire6(83);
	sub_wire2(0, 84)    <= sub_wire6(84);
	sub_wire2(0, 85)    <= sub_wire6(85);
	sub_wire2(0, 86)    <= sub_wire6(86);
	sub_wire2(0, 87)    <= sub_wire6(87);
	sub_wire2(0, 88)    <= sub_wire6(88);
	sub_wire2(0, 89)    <= sub_wire6(89);
	sub_wire2(0, 90)    <= sub_wire6(90);
	sub_wire2(0, 91)    <= sub_wire6(91);
	sub_wire2(0, 92)    <= sub_wire6(92);
	sub_wire2(0, 93)    <= sub_wire6(93);
	sub_wire2(0, 94)    <= sub_wire6(94);
	sub_wire2(0, 95)    <= sub_wire6(95);
	sub_wire2(0, 96)    <= sub_wire6(96);
	sub_wire2(0, 97)    <= sub_wire6(97);
	sub_wire2(0, 98)    <= sub_wire6(98);
	sub_wire2(0, 99)    <= sub_wire6(99);
	sub_wire2(0, 100)    <= sub_wire6(100);
	sub_wire2(0, 101)    <= sub_wire6(101);
	sub_wire2(0, 102)    <= sub_wire6(102);
	sub_wire2(0, 103)    <= sub_wire6(103);
	sub_wire2(0, 104)    <= sub_wire6(104);
	sub_wire2(0, 105)    <= sub_wire6(105);
	sub_wire2(0, 106)    <= sub_wire6(106);
	sub_wire2(0, 107)    <= sub_wire6(107);
	sub_wire2(0, 108)    <= sub_wire6(108);
	sub_wire2(0, 109)    <= sub_wire6(109);
	sub_wire2(0, 110)    <= sub_wire6(110);
	sub_wire2(0, 111)    <= sub_wire6(111);
	sub_wire2(0, 112)    <= sub_wire6(112);
	sub_wire2(0, 113)    <= sub_wire6(113);
	sub_wire2(0, 114)    <= sub_wire6(114);
	sub_wire2(0, 115)    <= sub_wire6(115);
	sub_wire2(0, 116)    <= sub_wire6(116);
	sub_wire2(0, 117)    <= sub_wire6(117);
	sub_wire2(0, 118)    <= sub_wire6(118);
	sub_wire2(0, 119)    <= sub_wire6(119);
	sub_wire2(0, 120)    <= sub_wire6(120);
	sub_wire2(0, 121)    <= sub_wire6(121);
	sub_wire2(0, 122)    <= sub_wire6(122);
	sub_wire2(0, 123)    <= sub_wire6(123);
	sub_wire2(0, 124)    <= sub_wire6(124);
	sub_wire2(0, 125)    <= sub_wire6(125);
	sub_wire2(0, 126)    <= sub_wire6(126);
	sub_wire2(0, 127)    <= sub_wire6(127);
	sub_wire2(0, 128)    <= sub_wire6(128);
	sub_wire2(0, 129)    <= sub_wire6(129);
	sub_wire2(0, 130)    <= sub_wire6(130);
	sub_wire2(0, 131)    <= sub_wire6(131);
	sub_wire2(0, 132)    <= sub_wire6(132);
	sub_wire2(0, 133)    <= sub_wire6(133);
	sub_wire2(0, 134)    <= sub_wire6(134);
	sub_wire2(0, 135)    <= sub_wire6(135);
	sub_wire2(0, 136)    <= sub_wire6(136);
	sub_wire2(0, 137)    <= sub_wire6(137);
	sub_wire2(0, 138)    <= sub_wire6(138);
	sub_wire2(0, 139)    <= sub_wire6(139);
	sub_wire2(0, 140)    <= sub_wire6(140);
	sub_wire2(0, 141)    <= sub_wire6(141);
	sub_wire2(0, 142)    <= sub_wire6(142);
	sub_wire2(0, 143)    <= sub_wire6(143);
	sub_wire2(0, 144)    <= sub_wire6(144);
	sub_wire2(0, 145)    <= sub_wire6(145);
	sub_wire2(0, 146)    <= sub_wire6(146);
	sub_wire2(0, 147)    <= sub_wire6(147);
	sub_wire2(0, 148)    <= sub_wire6(148);
	sub_wire2(0, 149)    <= sub_wire6(149);
	sub_wire2(0, 150)    <= sub_wire6(150);
	sub_wire2(0, 151)    <= sub_wire6(151);
	sub_wire2(0, 152)    <= sub_wire6(152);
	sub_wire2(0, 153)    <= sub_wire6(153);
	sub_wire2(0, 154)    <= sub_wire6(154);
	sub_wire2(0, 155)    <= sub_wire6(155);
	sub_wire2(0, 156)    <= sub_wire6(156);
	sub_wire2(0, 157)    <= sub_wire6(157);
	sub_wire2(0, 158)    <= sub_wire6(158);
	sub_wire2(0, 159)    <= sub_wire6(159);
	sub_wire2(0, 160)    <= sub_wire6(160);
	sub_wire2(0, 161)    <= sub_wire6(161);
	sub_wire2(0, 162)    <= sub_wire6(162);
	sub_wire2(0, 163)    <= sub_wire6(163);
	sub_wire2(0, 164)    <= sub_wire6(164);
	sub_wire2(0, 165)    <= sub_wire6(165);
	sub_wire2(0, 166)    <= sub_wire6(166);
	sub_wire2(0, 167)    <= sub_wire6(167);
	sub_wire2(0, 168)    <= sub_wire6(168);
	sub_wire2(0, 169)    <= sub_wire6(169);
	sub_wire2(0, 170)    <= sub_wire6(170);
	sub_wire2(0, 171)    <= sub_wire6(171);
	sub_wire2(0, 172)    <= sub_wire6(172);
	sub_wire2(0, 173)    <= sub_wire6(173);
	sub_wire2(0, 174)    <= sub_wire6(174);
	sub_wire2(0, 175)    <= sub_wire6(175);
	sub_wire2(0, 176)    <= sub_wire6(176);
	sub_wire2(0, 177)    <= sub_wire6(177);
	sub_wire2(0, 178)    <= sub_wire6(178);
	sub_wire2(0, 179)    <= sub_wire6(179);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_pipeline => 1,
		lpm_size => 5,
		lpm_type => "LPM_MUX",
		lpm_width => 180,
		lpm_widths => 3
	)
	PORT MAP (
		sel => sel,
		aclr => aclr,
		clock => clock,
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "5"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "180"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND aclr
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
-- Retrieval info: USED_PORT: data0x 0 0 180 0 INPUT NODEFVAL data0x[179..0]
-- Retrieval info: USED_PORT: data1x 0 0 180 0 INPUT NODEFVAL data1x[179..0]
-- Retrieval info: USED_PORT: data2x 0 0 180 0 INPUT NODEFVAL data2x[179..0]
-- Retrieval info: USED_PORT: data3x 0 0 180 0 INPUT NODEFVAL data3x[179..0]
-- Retrieval info: USED_PORT: data4x 0 0 180 0 INPUT NODEFVAL data4x[179..0]
-- Retrieval info: USED_PORT: result 0 0 180 0 OUTPUT NODEFVAL result[179..0]
-- Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL sel[2..0]
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 180 0 @result 0 0 180 0
-- Retrieval info: CONNECT: @data 1 4 180 0 data4x 0 0 180 0
-- Retrieval info: CONNECT: @data 1 3 180 0 data3x 0 0 180 0
-- Retrieval info: CONNECT: @data 1 2 180 0 data2x 0 0 180 0
-- Retrieval info: CONNECT: @data 1 1 180 0 data1x 0 0 180 0
-- Retrieval info: CONNECT: @data 1 0 180 0 data0x 0 0 180 0
-- Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_51_180_p1.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_51_180_p1.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_51_180_p1.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_51_180_p1.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_51_180_p1_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
