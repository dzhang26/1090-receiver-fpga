-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: mux_21_180.vhd
-- Megafunction Name(s):
-- 			lpm_mux
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux_21_180 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (179 DOWNTO 0);
		sel		: IN STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (179 DOWNTO 0)
	);
END mux_21_180;


ARCHITECTURE SYN OF mux_21_180 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (179 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_2D (1 DOWNTO 0, 179 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (179 DOWNTO 0);

BEGIN
	sub_wire5    <= data0x(179 DOWNTO 0);
	result    <= sub_wire0(179 DOWNTO 0);
	sub_wire1    <= sel;
	sub_wire2(0)    <= sub_wire1;
	sub_wire3    <= data1x(179 DOWNTO 0);
	sub_wire4(1, 0)    <= sub_wire3(0);
	sub_wire4(1, 1)    <= sub_wire3(1);
	sub_wire4(1, 2)    <= sub_wire3(2);
	sub_wire4(1, 3)    <= sub_wire3(3);
	sub_wire4(1, 4)    <= sub_wire3(4);
	sub_wire4(1, 5)    <= sub_wire3(5);
	sub_wire4(1, 6)    <= sub_wire3(6);
	sub_wire4(1, 7)    <= sub_wire3(7);
	sub_wire4(1, 8)    <= sub_wire3(8);
	sub_wire4(1, 9)    <= sub_wire3(9);
	sub_wire4(1, 10)    <= sub_wire3(10);
	sub_wire4(1, 11)    <= sub_wire3(11);
	sub_wire4(1, 12)    <= sub_wire3(12);
	sub_wire4(1, 13)    <= sub_wire3(13);
	sub_wire4(1, 14)    <= sub_wire3(14);
	sub_wire4(1, 15)    <= sub_wire3(15);
	sub_wire4(1, 16)    <= sub_wire3(16);
	sub_wire4(1, 17)    <= sub_wire3(17);
	sub_wire4(1, 18)    <= sub_wire3(18);
	sub_wire4(1, 19)    <= sub_wire3(19);
	sub_wire4(1, 20)    <= sub_wire3(20);
	sub_wire4(1, 21)    <= sub_wire3(21);
	sub_wire4(1, 22)    <= sub_wire3(22);
	sub_wire4(1, 23)    <= sub_wire3(23);
	sub_wire4(1, 24)    <= sub_wire3(24);
	sub_wire4(1, 25)    <= sub_wire3(25);
	sub_wire4(1, 26)    <= sub_wire3(26);
	sub_wire4(1, 27)    <= sub_wire3(27);
	sub_wire4(1, 28)    <= sub_wire3(28);
	sub_wire4(1, 29)    <= sub_wire3(29);
	sub_wire4(1, 30)    <= sub_wire3(30);
	sub_wire4(1, 31)    <= sub_wire3(31);
	sub_wire4(1, 32)    <= sub_wire3(32);
	sub_wire4(1, 33)    <= sub_wire3(33);
	sub_wire4(1, 34)    <= sub_wire3(34);
	sub_wire4(1, 35)    <= sub_wire3(35);
	sub_wire4(1, 36)    <= sub_wire3(36);
	sub_wire4(1, 37)    <= sub_wire3(37);
	sub_wire4(1, 38)    <= sub_wire3(38);
	sub_wire4(1, 39)    <= sub_wire3(39);
	sub_wire4(1, 40)    <= sub_wire3(40);
	sub_wire4(1, 41)    <= sub_wire3(41);
	sub_wire4(1, 42)    <= sub_wire3(42);
	sub_wire4(1, 43)    <= sub_wire3(43);
	sub_wire4(1, 44)    <= sub_wire3(44);
	sub_wire4(1, 45)    <= sub_wire3(45);
	sub_wire4(1, 46)    <= sub_wire3(46);
	sub_wire4(1, 47)    <= sub_wire3(47);
	sub_wire4(1, 48)    <= sub_wire3(48);
	sub_wire4(1, 49)    <= sub_wire3(49);
	sub_wire4(1, 50)    <= sub_wire3(50);
	sub_wire4(1, 51)    <= sub_wire3(51);
	sub_wire4(1, 52)    <= sub_wire3(52);
	sub_wire4(1, 53)    <= sub_wire3(53);
	sub_wire4(1, 54)    <= sub_wire3(54);
	sub_wire4(1, 55)    <= sub_wire3(55);
	sub_wire4(1, 56)    <= sub_wire3(56);
	sub_wire4(1, 57)    <= sub_wire3(57);
	sub_wire4(1, 58)    <= sub_wire3(58);
	sub_wire4(1, 59)    <= sub_wire3(59);
	sub_wire4(1, 60)    <= sub_wire3(60);
	sub_wire4(1, 61)    <= sub_wire3(61);
	sub_wire4(1, 62)    <= sub_wire3(62);
	sub_wire4(1, 63)    <= sub_wire3(63);
	sub_wire4(1, 64)    <= sub_wire3(64);
	sub_wire4(1, 65)    <= sub_wire3(65);
	sub_wire4(1, 66)    <= sub_wire3(66);
	sub_wire4(1, 67)    <= sub_wire3(67);
	sub_wire4(1, 68)    <= sub_wire3(68);
	sub_wire4(1, 69)    <= sub_wire3(69);
	sub_wire4(1, 70)    <= sub_wire3(70);
	sub_wire4(1, 71)    <= sub_wire3(71);
	sub_wire4(1, 72)    <= sub_wire3(72);
	sub_wire4(1, 73)    <= sub_wire3(73);
	sub_wire4(1, 74)    <= sub_wire3(74);
	sub_wire4(1, 75)    <= sub_wire3(75);
	sub_wire4(1, 76)    <= sub_wire3(76);
	sub_wire4(1, 77)    <= sub_wire3(77);
	sub_wire4(1, 78)    <= sub_wire3(78);
	sub_wire4(1, 79)    <= sub_wire3(79);
	sub_wire4(1, 80)    <= sub_wire3(80);
	sub_wire4(1, 81)    <= sub_wire3(81);
	sub_wire4(1, 82)    <= sub_wire3(82);
	sub_wire4(1, 83)    <= sub_wire3(83);
	sub_wire4(1, 84)    <= sub_wire3(84);
	sub_wire4(1, 85)    <= sub_wire3(85);
	sub_wire4(1, 86)    <= sub_wire3(86);
	sub_wire4(1, 87)    <= sub_wire3(87);
	sub_wire4(1, 88)    <= sub_wire3(88);
	sub_wire4(1, 89)    <= sub_wire3(89);
	sub_wire4(1, 90)    <= sub_wire3(90);
	sub_wire4(1, 91)    <= sub_wire3(91);
	sub_wire4(1, 92)    <= sub_wire3(92);
	sub_wire4(1, 93)    <= sub_wire3(93);
	sub_wire4(1, 94)    <= sub_wire3(94);
	sub_wire4(1, 95)    <= sub_wire3(95);
	sub_wire4(1, 96)    <= sub_wire3(96);
	sub_wire4(1, 97)    <= sub_wire3(97);
	sub_wire4(1, 98)    <= sub_wire3(98);
	sub_wire4(1, 99)    <= sub_wire3(99);
	sub_wire4(1, 100)    <= sub_wire3(100);
	sub_wire4(1, 101)    <= sub_wire3(101);
	sub_wire4(1, 102)    <= sub_wire3(102);
	sub_wire4(1, 103)    <= sub_wire3(103);
	sub_wire4(1, 104)    <= sub_wire3(104);
	sub_wire4(1, 105)    <= sub_wire3(105);
	sub_wire4(1, 106)    <= sub_wire3(106);
	sub_wire4(1, 107)    <= sub_wire3(107);
	sub_wire4(1, 108)    <= sub_wire3(108);
	sub_wire4(1, 109)    <= sub_wire3(109);
	sub_wire4(1, 110)    <= sub_wire3(110);
	sub_wire4(1, 111)    <= sub_wire3(111);
	sub_wire4(1, 112)    <= sub_wire3(112);
	sub_wire4(1, 113)    <= sub_wire3(113);
	sub_wire4(1, 114)    <= sub_wire3(114);
	sub_wire4(1, 115)    <= sub_wire3(115);
	sub_wire4(1, 116)    <= sub_wire3(116);
	sub_wire4(1, 117)    <= sub_wire3(117);
	sub_wire4(1, 118)    <= sub_wire3(118);
	sub_wire4(1, 119)    <= sub_wire3(119);
	sub_wire4(1, 120)    <= sub_wire3(120);
	sub_wire4(1, 121)    <= sub_wire3(121);
	sub_wire4(1, 122)    <= sub_wire3(122);
	sub_wire4(1, 123)    <= sub_wire3(123);
	sub_wire4(1, 124)    <= sub_wire3(124);
	sub_wire4(1, 125)    <= sub_wire3(125);
	sub_wire4(1, 126)    <= sub_wire3(126);
	sub_wire4(1, 127)    <= sub_wire3(127);
	sub_wire4(1, 128)    <= sub_wire3(128);
	sub_wire4(1, 129)    <= sub_wire3(129);
	sub_wire4(1, 130)    <= sub_wire3(130);
	sub_wire4(1, 131)    <= sub_wire3(131);
	sub_wire4(1, 132)    <= sub_wire3(132);
	sub_wire4(1, 133)    <= sub_wire3(133);
	sub_wire4(1, 134)    <= sub_wire3(134);
	sub_wire4(1, 135)    <= sub_wire3(135);
	sub_wire4(1, 136)    <= sub_wire3(136);
	sub_wire4(1, 137)    <= sub_wire3(137);
	sub_wire4(1, 138)    <= sub_wire3(138);
	sub_wire4(1, 139)    <= sub_wire3(139);
	sub_wire4(1, 140)    <= sub_wire3(140);
	sub_wire4(1, 141)    <= sub_wire3(141);
	sub_wire4(1, 142)    <= sub_wire3(142);
	sub_wire4(1, 143)    <= sub_wire3(143);
	sub_wire4(1, 144)    <= sub_wire3(144);
	sub_wire4(1, 145)    <= sub_wire3(145);
	sub_wire4(1, 146)    <= sub_wire3(146);
	sub_wire4(1, 147)    <= sub_wire3(147);
	sub_wire4(1, 148)    <= sub_wire3(148);
	sub_wire4(1, 149)    <= sub_wire3(149);
	sub_wire4(1, 150)    <= sub_wire3(150);
	sub_wire4(1, 151)    <= sub_wire3(151);
	sub_wire4(1, 152)    <= sub_wire3(152);
	sub_wire4(1, 153)    <= sub_wire3(153);
	sub_wire4(1, 154)    <= sub_wire3(154);
	sub_wire4(1, 155)    <= sub_wire3(155);
	sub_wire4(1, 156)    <= sub_wire3(156);
	sub_wire4(1, 157)    <= sub_wire3(157);
	sub_wire4(1, 158)    <= sub_wire3(158);
	sub_wire4(1, 159)    <= sub_wire3(159);
	sub_wire4(1, 160)    <= sub_wire3(160);
	sub_wire4(1, 161)    <= sub_wire3(161);
	sub_wire4(1, 162)    <= sub_wire3(162);
	sub_wire4(1, 163)    <= sub_wire3(163);
	sub_wire4(1, 164)    <= sub_wire3(164);
	sub_wire4(1, 165)    <= sub_wire3(165);
	sub_wire4(1, 166)    <= sub_wire3(166);
	sub_wire4(1, 167)    <= sub_wire3(167);
	sub_wire4(1, 168)    <= sub_wire3(168);
	sub_wire4(1, 169)    <= sub_wire3(169);
	sub_wire4(1, 170)    <= sub_wire3(170);
	sub_wire4(1, 171)    <= sub_wire3(171);
	sub_wire4(1, 172)    <= sub_wire3(172);
	sub_wire4(1, 173)    <= sub_wire3(173);
	sub_wire4(1, 174)    <= sub_wire3(174);
	sub_wire4(1, 175)    <= sub_wire3(175);
	sub_wire4(1, 176)    <= sub_wire3(176);
	sub_wire4(1, 177)    <= sub_wire3(177);
	sub_wire4(1, 178)    <= sub_wire3(178);
	sub_wire4(1, 179)    <= sub_wire3(179);
	sub_wire4(0, 0)    <= sub_wire5(0);
	sub_wire4(0, 1)    <= sub_wire5(1);
	sub_wire4(0, 2)    <= sub_wire5(2);
	sub_wire4(0, 3)    <= sub_wire5(3);
	sub_wire4(0, 4)    <= sub_wire5(4);
	sub_wire4(0, 5)    <= sub_wire5(5);
	sub_wire4(0, 6)    <= sub_wire5(6);
	sub_wire4(0, 7)    <= sub_wire5(7);
	sub_wire4(0, 8)    <= sub_wire5(8);
	sub_wire4(0, 9)    <= sub_wire5(9);
	sub_wire4(0, 10)    <= sub_wire5(10);
	sub_wire4(0, 11)    <= sub_wire5(11);
	sub_wire4(0, 12)    <= sub_wire5(12);
	sub_wire4(0, 13)    <= sub_wire5(13);
	sub_wire4(0, 14)    <= sub_wire5(14);
	sub_wire4(0, 15)    <= sub_wire5(15);
	sub_wire4(0, 16)    <= sub_wire5(16);
	sub_wire4(0, 17)    <= sub_wire5(17);
	sub_wire4(0, 18)    <= sub_wire5(18);
	sub_wire4(0, 19)    <= sub_wire5(19);
	sub_wire4(0, 20)    <= sub_wire5(20);
	sub_wire4(0, 21)    <= sub_wire5(21);
	sub_wire4(0, 22)    <= sub_wire5(22);
	sub_wire4(0, 23)    <= sub_wire5(23);
	sub_wire4(0, 24)    <= sub_wire5(24);
	sub_wire4(0, 25)    <= sub_wire5(25);
	sub_wire4(0, 26)    <= sub_wire5(26);
	sub_wire4(0, 27)    <= sub_wire5(27);
	sub_wire4(0, 28)    <= sub_wire5(28);
	sub_wire4(0, 29)    <= sub_wire5(29);
	sub_wire4(0, 30)    <= sub_wire5(30);
	sub_wire4(0, 31)    <= sub_wire5(31);
	sub_wire4(0, 32)    <= sub_wire5(32);
	sub_wire4(0, 33)    <= sub_wire5(33);
	sub_wire4(0, 34)    <= sub_wire5(34);
	sub_wire4(0, 35)    <= sub_wire5(35);
	sub_wire4(0, 36)    <= sub_wire5(36);
	sub_wire4(0, 37)    <= sub_wire5(37);
	sub_wire4(0, 38)    <= sub_wire5(38);
	sub_wire4(0, 39)    <= sub_wire5(39);
	sub_wire4(0, 40)    <= sub_wire5(40);
	sub_wire4(0, 41)    <= sub_wire5(41);
	sub_wire4(0, 42)    <= sub_wire5(42);
	sub_wire4(0, 43)    <= sub_wire5(43);
	sub_wire4(0, 44)    <= sub_wire5(44);
	sub_wire4(0, 45)    <= sub_wire5(45);
	sub_wire4(0, 46)    <= sub_wire5(46);
	sub_wire4(0, 47)    <= sub_wire5(47);
	sub_wire4(0, 48)    <= sub_wire5(48);
	sub_wire4(0, 49)    <= sub_wire5(49);
	sub_wire4(0, 50)    <= sub_wire5(50);
	sub_wire4(0, 51)    <= sub_wire5(51);
	sub_wire4(0, 52)    <= sub_wire5(52);
	sub_wire4(0, 53)    <= sub_wire5(53);
	sub_wire4(0, 54)    <= sub_wire5(54);
	sub_wire4(0, 55)    <= sub_wire5(55);
	sub_wire4(0, 56)    <= sub_wire5(56);
	sub_wire4(0, 57)    <= sub_wire5(57);
	sub_wire4(0, 58)    <= sub_wire5(58);
	sub_wire4(0, 59)    <= sub_wire5(59);
	sub_wire4(0, 60)    <= sub_wire5(60);
	sub_wire4(0, 61)    <= sub_wire5(61);
	sub_wire4(0, 62)    <= sub_wire5(62);
	sub_wire4(0, 63)    <= sub_wire5(63);
	sub_wire4(0, 64)    <= sub_wire5(64);
	sub_wire4(0, 65)    <= sub_wire5(65);
	sub_wire4(0, 66)    <= sub_wire5(66);
	sub_wire4(0, 67)    <= sub_wire5(67);
	sub_wire4(0, 68)    <= sub_wire5(68);
	sub_wire4(0, 69)    <= sub_wire5(69);
	sub_wire4(0, 70)    <= sub_wire5(70);
	sub_wire4(0, 71)    <= sub_wire5(71);
	sub_wire4(0, 72)    <= sub_wire5(72);
	sub_wire4(0, 73)    <= sub_wire5(73);
	sub_wire4(0, 74)    <= sub_wire5(74);
	sub_wire4(0, 75)    <= sub_wire5(75);
	sub_wire4(0, 76)    <= sub_wire5(76);
	sub_wire4(0, 77)    <= sub_wire5(77);
	sub_wire4(0, 78)    <= sub_wire5(78);
	sub_wire4(0, 79)    <= sub_wire5(79);
	sub_wire4(0, 80)    <= sub_wire5(80);
	sub_wire4(0, 81)    <= sub_wire5(81);
	sub_wire4(0, 82)    <= sub_wire5(82);
	sub_wire4(0, 83)    <= sub_wire5(83);
	sub_wire4(0, 84)    <= sub_wire5(84);
	sub_wire4(0, 85)    <= sub_wire5(85);
	sub_wire4(0, 86)    <= sub_wire5(86);
	sub_wire4(0, 87)    <= sub_wire5(87);
	sub_wire4(0, 88)    <= sub_wire5(88);
	sub_wire4(0, 89)    <= sub_wire5(89);
	sub_wire4(0, 90)    <= sub_wire5(90);
	sub_wire4(0, 91)    <= sub_wire5(91);
	sub_wire4(0, 92)    <= sub_wire5(92);
	sub_wire4(0, 93)    <= sub_wire5(93);
	sub_wire4(0, 94)    <= sub_wire5(94);
	sub_wire4(0, 95)    <= sub_wire5(95);
	sub_wire4(0, 96)    <= sub_wire5(96);
	sub_wire4(0, 97)    <= sub_wire5(97);
	sub_wire4(0, 98)    <= sub_wire5(98);
	sub_wire4(0, 99)    <= sub_wire5(99);
	sub_wire4(0, 100)    <= sub_wire5(100);
	sub_wire4(0, 101)    <= sub_wire5(101);
	sub_wire4(0, 102)    <= sub_wire5(102);
	sub_wire4(0, 103)    <= sub_wire5(103);
	sub_wire4(0, 104)    <= sub_wire5(104);
	sub_wire4(0, 105)    <= sub_wire5(105);
	sub_wire4(0, 106)    <= sub_wire5(106);
	sub_wire4(0, 107)    <= sub_wire5(107);
	sub_wire4(0, 108)    <= sub_wire5(108);
	sub_wire4(0, 109)    <= sub_wire5(109);
	sub_wire4(0, 110)    <= sub_wire5(110);
	sub_wire4(0, 111)    <= sub_wire5(111);
	sub_wire4(0, 112)    <= sub_wire5(112);
	sub_wire4(0, 113)    <= sub_wire5(113);
	sub_wire4(0, 114)    <= sub_wire5(114);
	sub_wire4(0, 115)    <= sub_wire5(115);
	sub_wire4(0, 116)    <= sub_wire5(116);
	sub_wire4(0, 117)    <= sub_wire5(117);
	sub_wire4(0, 118)    <= sub_wire5(118);
	sub_wire4(0, 119)    <= sub_wire5(119);
	sub_wire4(0, 120)    <= sub_wire5(120);
	sub_wire4(0, 121)    <= sub_wire5(121);
	sub_wire4(0, 122)    <= sub_wire5(122);
	sub_wire4(0, 123)    <= sub_wire5(123);
	sub_wire4(0, 124)    <= sub_wire5(124);
	sub_wire4(0, 125)    <= sub_wire5(125);
	sub_wire4(0, 126)    <= sub_wire5(126);
	sub_wire4(0, 127)    <= sub_wire5(127);
	sub_wire4(0, 128)    <= sub_wire5(128);
	sub_wire4(0, 129)    <= sub_wire5(129);
	sub_wire4(0, 130)    <= sub_wire5(130);
	sub_wire4(0, 131)    <= sub_wire5(131);
	sub_wire4(0, 132)    <= sub_wire5(132);
	sub_wire4(0, 133)    <= sub_wire5(133);
	sub_wire4(0, 134)    <= sub_wire5(134);
	sub_wire4(0, 135)    <= sub_wire5(135);
	sub_wire4(0, 136)    <= sub_wire5(136);
	sub_wire4(0, 137)    <= sub_wire5(137);
	sub_wire4(0, 138)    <= sub_wire5(138);
	sub_wire4(0, 139)    <= sub_wire5(139);
	sub_wire4(0, 140)    <= sub_wire5(140);
	sub_wire4(0, 141)    <= sub_wire5(141);
	sub_wire4(0, 142)    <= sub_wire5(142);
	sub_wire4(0, 143)    <= sub_wire5(143);
	sub_wire4(0, 144)    <= sub_wire5(144);
	sub_wire4(0, 145)    <= sub_wire5(145);
	sub_wire4(0, 146)    <= sub_wire5(146);
	sub_wire4(0, 147)    <= sub_wire5(147);
	sub_wire4(0, 148)    <= sub_wire5(148);
	sub_wire4(0, 149)    <= sub_wire5(149);
	sub_wire4(0, 150)    <= sub_wire5(150);
	sub_wire4(0, 151)    <= sub_wire5(151);
	sub_wire4(0, 152)    <= sub_wire5(152);
	sub_wire4(0, 153)    <= sub_wire5(153);
	sub_wire4(0, 154)    <= sub_wire5(154);
	sub_wire4(0, 155)    <= sub_wire5(155);
	sub_wire4(0, 156)    <= sub_wire5(156);
	sub_wire4(0, 157)    <= sub_wire5(157);
	sub_wire4(0, 158)    <= sub_wire5(158);
	sub_wire4(0, 159)    <= sub_wire5(159);
	sub_wire4(0, 160)    <= sub_wire5(160);
	sub_wire4(0, 161)    <= sub_wire5(161);
	sub_wire4(0, 162)    <= sub_wire5(162);
	sub_wire4(0, 163)    <= sub_wire5(163);
	sub_wire4(0, 164)    <= sub_wire5(164);
	sub_wire4(0, 165)    <= sub_wire5(165);
	sub_wire4(0, 166)    <= sub_wire5(166);
	sub_wire4(0, 167)    <= sub_wire5(167);
	sub_wire4(0, 168)    <= sub_wire5(168);
	sub_wire4(0, 169)    <= sub_wire5(169);
	sub_wire4(0, 170)    <= sub_wire5(170);
	sub_wire4(0, 171)    <= sub_wire5(171);
	sub_wire4(0, 172)    <= sub_wire5(172);
	sub_wire4(0, 173)    <= sub_wire5(173);
	sub_wire4(0, 174)    <= sub_wire5(174);
	sub_wire4(0, 175)    <= sub_wire5(175);
	sub_wire4(0, 176)    <= sub_wire5(176);
	sub_wire4(0, 177)    <= sub_wire5(177);
	sub_wire4(0, 178)    <= sub_wire5(178);
	sub_wire4(0, 179)    <= sub_wire5(179);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_size => 2,
		lpm_type => "LPM_MUX",
		lpm_width => 180,
		lpm_widths => 1
	)
	PORT MAP (
		sel => sub_wire2,
		data => sub_wire4,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "180"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
-- Retrieval info: USED_PORT: data0x 0 0 180 0 INPUT NODEFVAL data0x[179..0]
-- Retrieval info: USED_PORT: data1x 0 0 180 0 INPUT NODEFVAL data1x[179..0]
-- Retrieval info: USED_PORT: result 0 0 180 0 OUTPUT NODEFVAL result[179..0]
-- Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL sel
-- Retrieval info: CONNECT: result 0 0 180 0 @result 0 0 180 0
-- Retrieval info: CONNECT: @data 1 1 180 0 data1x 0 0 180 0
-- Retrieval info: CONNECT: @data 1 0 180 0 data0x 0 0 180 0
-- Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_21_180.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_21_180.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_21_180.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_21_180.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux_21_180_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
